<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-51.5371,-510.455,40.2629,-555.83</PageViewport>
<gate>
<ID>390</ID>
<type>GA_LED</type>
<position>-9,-541.5</position>
<input>
<ID>N_in0</ID>154 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2</ID>
<type>AA_MUX_2x1</type>
<position>34.5,-12.5</position>
<input>
<ID>IN_0</ID>3 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>5 </output>
<input>
<ID>SEL_0</ID>4 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>392</ID>
<type>GA_LED</type>
<position>-9,-549</position>
<input>
<ID>N_in0</ID>155 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>394</ID>
<type>AI_XOR2</type>
<position>-24.5,-540.5</position>
<input>
<ID>IN_0</ID>152 </input>
<input>
<ID>IN_1</ID>156 </input>
<output>
<ID>OUT</ID>154 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6</ID>
<type>AA_TOGGLE</type>
<position>16,-10.5</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>396</ID>
<type>AI_XOR2</type>
<position>-17,-549</position>
<input>
<ID>IN_0</ID>154 </input>
<input>
<ID>IN_1</ID>153 </input>
<output>
<ID>OUT</ID>155 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>8</ID>
<type>AA_TOGGLE</type>
<position>16,-17</position>
<output>
<ID>OUT_0</ID>3 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>10</ID>
<type>AA_TOGGLE</type>
<position>34.5,-5</position>
<output>
<ID>OUT_0</ID>4 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>12</ID>
<type>GA_LED</type>
<position>37.5,-12.5</position>
<input>
<ID>N_in0</ID>5 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>14</ID>
<type>AE_MUX_4x1</type>
<position>83,-14.5</position>
<input>
<ID>IN_0</ID>9 </input>
<input>
<ID>IN_1</ID>8 </input>
<input>
<ID>IN_2</ID>7 </input>
<input>
<ID>IN_3</ID>6 </input>
<output>
<ID>OUT</ID>12 </output>
<input>
<ID>SEL_0</ID>11 </input>
<input>
<ID>SEL_1</ID>10 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>16</ID>
<type>AA_TOGGLE</type>
<position>67,-9.5</position>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>18</ID>
<type>AA_TOGGLE</type>
<position>67,-13.5</position>
<output>
<ID>OUT_0</ID>7 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>20</ID>
<type>AA_TOGGLE</type>
<position>61,-16</position>
<output>
<ID>OUT_0</ID>8 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>22</ID>
<type>AA_TOGGLE</type>
<position>67,-19.5</position>
<output>
<ID>OUT_0</ID>9 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>24</ID>
<type>AA_TOGGLE</type>
<position>83,-4.5</position>
<output>
<ID>OUT_0</ID>10 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>26</ID>
<type>AA_TOGGLE</type>
<position>90,-3.5</position>
<output>
<ID>OUT_0</ID>11 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>28</ID>
<type>GA_LED</type>
<position>100.5,-14.5</position>
<input>
<ID>N_in0</ID>12 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>30</ID>
<type>AI_MUX_8x1</type>
<position>35,-42</position>
<input>
<ID>IN_0</ID>19 </input>
<input>
<ID>IN_1</ID>18 </input>
<input>
<ID>IN_2</ID>17 </input>
<input>
<ID>IN_4</ID>16 </input>
<input>
<ID>IN_5</ID>15 </input>
<input>
<ID>IN_6</ID>14 </input>
<input>
<ID>IN_7</ID>13 </input>
<output>
<ID>OUT</ID>23 </output>
<input>
<ID>SEL_0</ID>22 </input>
<input>
<ID>SEL_1</ID>21 </input>
<input>
<ID>SEL_2</ID>20 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>32</ID>
<type>AA_TOGGLE</type>
<position>23.5,-32.5</position>
<output>
<ID>OUT_0</ID>13 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>34</ID>
<type>AA_TOGGLE</type>
<position>23.5,-39.5</position>
<output>
<ID>OUT_0</ID>14 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>36</ID>
<type>AA_TOGGLE</type>
<position>23.5,-36</position>
<output>
<ID>OUT_0</ID>15 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>38</ID>
<type>AA_TOGGLE</type>
<position>23,-42.5</position>
<output>
<ID>OUT_0</ID>16 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>40</ID>
<type>AA_TOGGLE</type>
<position>17,-44</position>
<output>
<ID>OUT_0</ID>17 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>42</ID>
<type>AA_TOGGLE</type>
<position>21.5,-47.5</position>
<output>
<ID>OUT_0</ID>18 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>44</ID>
<type>AA_TOGGLE</type>
<position>27.5,-50</position>
<output>
<ID>OUT_0</ID>19 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>46</ID>
<type>AA_TOGGLE</type>
<position>32.5,-28.5</position>
<output>
<ID>OUT_0</ID>20 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>48</ID>
<type>AA_TOGGLE</type>
<position>35,-28.5</position>
<output>
<ID>OUT_0</ID>21 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>50</ID>
<type>AA_TOGGLE</type>
<position>38.5,-28.5</position>
<output>
<ID>OUT_0</ID>22 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>52</ID>
<type>GA_LED</type>
<position>39,-42</position>
<input>
<ID>N_in0</ID>23 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>54</ID>
<type>AA_LABEL</type>
<position>10,-3</position>
<gparam>LABEL_TEXT 2x1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>56</ID>
<type>AA_LABEL</type>
<position>104,-5.5</position>
<gparam>LABEL_TEXT 4x1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>58</ID>
<type>AA_LABEL</type>
<position>28,-26</position>
<gparam>LABEL_TEXT 8x1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>60</ID>
<type>AA_LABEL</type>
<position>10,-10</position>
<gparam>LABEL_TEXT D1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>61</ID>
<type>AA_LABEL</type>
<position>11,-17</position>
<gparam>LABEL_TEXT D0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>62</ID>
<type>AA_LABEL</type>
<position>63,-10</position>
<gparam>LABEL_TEXT D3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>63</ID>
<type>AA_LABEL</type>
<position>63.5,-13.5</position>
<gparam>LABEL_TEXT D2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>64</ID>
<type>AA_LABEL</type>
<position>63.5,-19</position>
<gparam>LABEL_TEXT D0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>65</ID>
<type>AA_LABEL</type>
<position>58,-16</position>
<gparam>LABEL_TEXT D1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>66</ID>
<type>AA_LABEL</type>
<position>24,-50</position>
<gparam>LABEL_TEXT D0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>67</ID>
<type>AA_LABEL</type>
<position>18,-47</position>
<gparam>LABEL_TEXT D1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>68</ID>
<type>AA_LABEL</type>
<position>14,-43.5</position>
<gparam>LABEL_TEXT D2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>69</ID>
<type>AA_LABEL</type>
<position>20.5,-42.5</position>
<gparam>LABEL_TEXT D3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>70</ID>
<type>AA_LABEL</type>
<position>20.5,-39</position>
<gparam>LABEL_TEXT D4</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>71</ID>
<type>AA_LABEL</type>
<position>20.5,-36</position>
<gparam>LABEL_TEXT D5</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>72</ID>
<type>AA_LABEL</type>
<position>20,-32.5</position>
<gparam>LABEL_TEXT D6</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>74</ID>
<type>AA_MUX_2x1</type>
<position>11.5,-64.5</position>
<input>
<ID>IN_0</ID>25 </input>
<input>
<ID>IN_1</ID>24 </input>
<output>
<ID>OUT</ID>40 </output>
<input>
<ID>SEL_0</ID>33 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>76</ID>
<type>AA_MUX_2x1</type>
<position>11.5,-73</position>
<input>
<ID>IN_0</ID>27 </input>
<input>
<ID>IN_1</ID>26 </input>
<output>
<ID>OUT</ID>41 </output>
<input>
<ID>SEL_0</ID>33 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>78</ID>
<type>AA_MUX_2x1</type>
<position>11.5,-81.5</position>
<input>
<ID>IN_0</ID>29 </input>
<input>
<ID>IN_1</ID>28 </input>
<output>
<ID>OUT</ID>42 </output>
<input>
<ID>SEL_0</ID>33 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>80</ID>
<type>AA_MUX_2x1</type>
<position>11.5,-91</position>
<input>
<ID>IN_0</ID>31 </input>
<input>
<ID>IN_1</ID>30 </input>
<output>
<ID>OUT</ID>43 </output>
<input>
<ID>SEL_0</ID>33 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>82</ID>
<type>AA_TOGGLE</type>
<position>1.5,-62.5</position>
<output>
<ID>OUT_0</ID>24 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>84</ID>
<type>AA_TOGGLE</type>
<position>2,-66</position>
<output>
<ID>OUT_0</ID>25 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>86</ID>
<type>AA_TOGGLE</type>
<position>2,-71</position>
<output>
<ID>OUT_0</ID>26 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>88</ID>
<type>AA_TOGGLE</type>
<position>2,-74.5</position>
<output>
<ID>OUT_0</ID>27 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>90</ID>
<type>AA_TOGGLE</type>
<position>2.5,-80</position>
<output>
<ID>OUT_0</ID>28 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>92</ID>
<type>AA_TOGGLE</type>
<position>2.5,-82.5</position>
<output>
<ID>OUT_0</ID>29 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>94</ID>
<type>AA_TOGGLE</type>
<position>3,-89</position>
<output>
<ID>OUT_0</ID>30 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>96</ID>
<type>AA_TOGGLE</type>
<position>3,-92.5</position>
<output>
<ID>OUT_0</ID>31 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>98</ID>
<type>AA_TOGGLE</type>
<position>13.5,-56.5</position>
<output>
<ID>OUT_0</ID>33 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>100</ID>
<type>AA_MUX_2x1</type>
<position>41.5,-65.5</position>
<input>
<ID>IN_0</ID>41 </input>
<input>
<ID>IN_1</ID>40 </input>
<output>
<ID>OUT</ID>45 </output>
<input>
<ID>SEL_0</ID>38 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>102</ID>
<type>AA_MUX_2x1</type>
<position>43,-78.5</position>
<input>
<ID>IN_0</ID>43 </input>
<input>
<ID>IN_1</ID>42 </input>
<output>
<ID>OUT</ID>44 </output>
<input>
<ID>SEL_0</ID>38 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>112</ID>
<type>AA_TOGGLE</type>
<position>43.5,-57.5</position>
<output>
<ID>OUT_0</ID>38 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>116</ID>
<type>AA_MUX_2x1</type>
<position>59.5,-72</position>
<input>
<ID>IN_0</ID>44 </input>
<input>
<ID>IN_1</ID>45 </input>
<output>
<ID>OUT</ID>46 </output>
<input>
<ID>SEL_0</ID>39 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>118</ID>
<type>AA_TOGGLE</type>
<position>59.5,-57.5</position>
<output>
<ID>OUT_0</ID>39 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>120</ID>
<type>GA_LED</type>
<position>62.5,-72</position>
<input>
<ID>N_in0</ID>46 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>121</ID>
<type>AA_LABEL</type>
<position>-1,-92.5</position>
<gparam>LABEL_TEXT D0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>122</ID>
<type>AA_LABEL</type>
<position>-1.5,-89</position>
<gparam>LABEL_TEXT D1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>123</ID>
<type>AA_LABEL</type>
<position>-1,-82.5</position>
<gparam>LABEL_TEXT D2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>124</ID>
<type>AA_LABEL</type>
<position>-2,-79.5</position>
<gparam>LABEL_TEXT D3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>125</ID>
<type>AA_LABEL</type>
<position>-2,-74.5</position>
<gparam>LABEL_TEXT D4</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>126</ID>
<type>AA_LABEL</type>
<position>-2,-71</position>
<gparam>LABEL_TEXT D5</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>127</ID>
<type>AA_LABEL</type>
<position>-2.5,-66</position>
<gparam>LABEL_TEXT D6</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>128</ID>
<type>AA_LABEL</type>
<position>-3,-62</position>
<gparam>LABEL_TEXT D7</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>130</ID>
<type>AA_TOGGLE</type>
<position>-16,-99.5</position>
<output>
<ID>OUT_0</ID>57 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>132</ID>
<type>AA_TOGGLE</type>
<position>5,-99.5</position>
<output>
<ID>OUT_0</ID>48 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>134</ID>
<type>AA_TOGGLE</type>
<position>23.5,-100.5</position>
<output>
<ID>OUT_0</ID>52 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>136</ID>
<type>AE_SMALL_INVERTER</type>
<position>-12,-105</position>
<input>
<ID>IN_0</ID>57 </input>
<output>
<ID>OUT_0</ID>50 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>138</ID>
<type>AE_SMALL_INVERTER</type>
<position>10,-104</position>
<input>
<ID>IN_0</ID>48 </input>
<output>
<ID>OUT_0</ID>58 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>148</ID>
<type>AA_AND3</type>
<position>43,-107</position>
<input>
<ID>IN_0</ID>52 </input>
<input>
<ID>IN_2</ID>50 </input>
<output>
<ID>OUT</ID>53 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>150</ID>
<type>AA_AND3</type>
<position>44,-120</position>
<input>
<ID>IN_0</ID>52 </input>
<input>
<ID>IN_1</ID>48 </input>
<input>
<ID>IN_2</ID>50 </input>
<output>
<ID>OUT</ID>54 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>152</ID>
<type>AA_AND3</type>
<position>43.5,-131.5</position>
<input>
<ID>IN_0</ID>52 </input>
<input>
<ID>IN_1</ID>58 </input>
<input>
<ID>IN_2</ID>57 </input>
<output>
<ID>OUT</ID>55 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>154</ID>
<type>AA_AND3</type>
<position>44.5,-143</position>
<input>
<ID>IN_0</ID>52 </input>
<input>
<ID>IN_1</ID>48 </input>
<input>
<ID>IN_2</ID>57 </input>
<output>
<ID>OUT</ID>56 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>155</ID>
<type>AA_LABEL</type>
<position>-16,-96.5</position>
<gparam>LABEL_TEXT s1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>156</ID>
<type>AA_LABEL</type>
<position>5.5,-97</position>
<gparam>LABEL_TEXT s0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>157</ID>
<type>AA_LABEL</type>
<position>23.5,-97.5</position>
<gparam>LABEL_TEXT Din</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>159</ID>
<type>GA_LED</type>
<position>47,-107</position>
<input>
<ID>N_in0</ID>53 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>161</ID>
<type>GA_LED</type>
<position>48,-120</position>
<input>
<ID>N_in0</ID>54 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>163</ID>
<type>GA_LED</type>
<position>47.5,-131.5</position>
<input>
<ID>N_in0</ID>55 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>165</ID>
<type>GA_LED</type>
<position>48.5,-143</position>
<input>
<ID>N_in0</ID>56 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>167</ID>
<type>AA_TOGGLE</type>
<position>-69,-168</position>
<output>
<ID>OUT_0</ID>69 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>169</ID>
<type>AA_TOGGLE</type>
<position>-52,-167.5</position>
<output>
<ID>OUT_0</ID>70 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>171</ID>
<type>AA_TOGGLE</type>
<position>-32.5,-167.5</position>
<output>
<ID>OUT_0</ID>71 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>173</ID>
<type>AA_TOGGLE</type>
<position>-11.5,-167.5</position>
<output>
<ID>OUT_0</ID>68 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>175</ID>
<type>AA_AND4</type>
<position>31,-173.5</position>
<input>
<ID>IN_0</ID>68 </input>
<input>
<ID>IN_1</ID>72 </input>
<input>
<ID>IN_2</ID>73 </input>
<input>
<ID>IN_3</ID>74 </input>
<output>
<ID>OUT</ID>82 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>177</ID>
<type>AA_AND4</type>
<position>41.5,-185</position>
<input>
<ID>IN_0</ID>68 </input>
<input>
<ID>IN_1</ID>71 </input>
<input>
<ID>IN_2</ID>73 </input>
<input>
<ID>IN_3</ID>74 </input>
<output>
<ID>OUT</ID>81 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>179</ID>
<type>AA_AND4</type>
<position>48.5,-196.5</position>
<input>
<ID>IN_0</ID>68 </input>
<input>
<ID>IN_1</ID>72 </input>
<input>
<ID>IN_2</ID>70 </input>
<input>
<ID>IN_3</ID>74 </input>
<output>
<ID>OUT</ID>80 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>181</ID>
<type>AA_AND4</type>
<position>51,-208.5</position>
<input>
<ID>IN_0</ID>68 </input>
<input>
<ID>IN_1</ID>70 </input>
<input>
<ID>IN_2</ID>71 </input>
<input>
<ID>IN_3</ID>74 </input>
<output>
<ID>OUT</ID>79 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>183</ID>
<type>AA_AND4</type>
<position>42,-223.5</position>
<input>
<ID>IN_0</ID>68 </input>
<input>
<ID>IN_1</ID>72 </input>
<input>
<ID>IN_2</ID>70 </input>
<input>
<ID>IN_3</ID>69 </input>
<output>
<ID>OUT</ID>78 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>185</ID>
<type>AA_AND4</type>
<position>47,-237.5</position>
<input>
<ID>IN_0</ID>68 </input>
<input>
<ID>IN_1</ID>71 </input>
<input>
<ID>IN_2</ID>69 </input>
<input>
<ID>IN_3</ID>69 </input>
<output>
<ID>OUT</ID>77 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>187</ID>
<type>AA_AND4</type>
<position>46,-250</position>
<input>
<ID>IN_0</ID>68 </input>
<input>
<ID>IN_1</ID>72 </input>
<input>
<ID>IN_2</ID>70 </input>
<input>
<ID>IN_3</ID>69 </input>
<output>
<ID>OUT</ID>76 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>189</ID>
<type>AA_AND4</type>
<position>48.5,-262</position>
<input>
<ID>IN_0</ID>68 </input>
<input>
<ID>IN_1</ID>69 </input>
<input>
<ID>IN_2</ID>70 </input>
<input>
<ID>IN_3</ID>71 </input>
<output>
<ID>OUT</ID>75 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>207</ID>
<type>AE_SMALL_INVERTER</type>
<position>-63.5,-172</position>
<input>
<ID>IN_0</ID>69 </input>
<output>
<ID>OUT_0</ID>74 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>209</ID>
<type>AE_SMALL_INVERTER</type>
<position>-46.5,-171</position>
<input>
<ID>IN_0</ID>70 </input>
<output>
<ID>OUT_0</ID>73 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>211</ID>
<type>AE_SMALL_INVERTER</type>
<position>-28,-170.5</position>
<input>
<ID>IN_0</ID>71 </input>
<output>
<ID>OUT_0</ID>72 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>212</ID>
<type>GA_LED</type>
<position>52.5,-262</position>
<input>
<ID>N_in0</ID>75 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>213</ID>
<type>GA_LED</type>
<position>50,-250</position>
<input>
<ID>N_in0</ID>76 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>214</ID>
<type>GA_LED</type>
<position>51,-237.5</position>
<input>
<ID>N_in0</ID>77 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>215</ID>
<type>GA_LED</type>
<position>46,-223.5</position>
<input>
<ID>N_in0</ID>78 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>216</ID>
<type>GA_LED</type>
<position>55,-208.5</position>
<input>
<ID>N_in0</ID>79 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>218</ID>
<type>GA_LED</type>
<position>52.5,-196.5</position>
<input>
<ID>N_in0</ID>80 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>219</ID>
<type>GA_LED</type>
<position>45.5,-185</position>
<input>
<ID>N_in0</ID>81 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>220</ID>
<type>GA_LED</type>
<position>35,-173.5</position>
<input>
<ID>N_in0</ID>82 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>222</ID>
<type>AA_TOGGLE</type>
<position>-94,-297</position>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>224</ID>
<type>AA_TOGGLE</type>
<position>-77.5,-297.5</position>
<output>
<ID>OUT_0</ID>90 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>226</ID>
<type>AA_TOGGLE</type>
<position>-64.5,-297</position>
<output>
<ID>OUT_0</ID>87 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>228</ID>
<type>AA_TOGGLE</type>
<position>-54.5,-297.5</position>
<output>
<ID>OUT_0</ID>88 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>230</ID>
<type>AA_TOGGLE</type>
<position>-43.5,-297.5</position>
<output>
<ID>OUT_0</ID>86 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>232</ID>
<type>AA_TOGGLE</type>
<position>-33,-297</position>
<output>
<ID>OUT_0</ID>85 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>234</ID>
<type>AA_TOGGLE</type>
<position>-23.5,-297</position>
<output>
<ID>OUT_0</ID>84 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>236</ID>
<type>AA_TOGGLE</type>
<position>-10.5,-297.5</position>
<output>
<ID>OUT_0</ID>83 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>238</ID>
<type>AE_OR4</type>
<position>32.5,-307</position>
<input>
<ID>IN_0</ID>83 </input>
<input>
<ID>IN_1</ID>84 </input>
<input>
<ID>IN_2</ID>85 </input>
<input>
<ID>IN_3</ID>86 </input>
<output>
<ID>OUT</ID>91 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>242</ID>
<type>AE_OR4</type>
<position>33,-337</position>
<input>
<ID>IN_0</ID>87 </input>
<input>
<ID>IN_1</ID>88 </input>
<input>
<ID>IN_2</ID>84 </input>
<input>
<ID>IN_3</ID>83 </input>
<output>
<ID>OUT</ID>92 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>244</ID>
<type>AE_OR4</type>
<position>34,-364.5</position>
<input>
<ID>IN_0</ID>90 </input>
<input>
<ID>IN_1</ID>88 </input>
<input>
<ID>IN_2</ID>85 </input>
<input>
<ID>IN_3</ID>83 </input>
<output>
<ID>OUT</ID>93 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>246</ID>
<type>GA_LED</type>
<position>37.5,-307</position>
<input>
<ID>N_in0</ID>91 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>248</ID>
<type>GA_LED</type>
<position>38,-337</position>
<input>
<ID>N_in0</ID>92 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>250</ID>
<type>GA_LED</type>
<position>39,-364.5</position>
<input>
<ID>N_in0</ID>93 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>252</ID>
<type>AA_TOGGLE</type>
<position>-85,-390</position>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>254</ID>
<type>AA_TOGGLE</type>
<position>-70,-390.5</position>
<output>
<ID>OUT_0</ID>98 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>256</ID>
<type>AA_TOGGLE</type>
<position>-56,-390.5</position>
<output>
<ID>OUT_0</ID>96 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>258</ID>
<type>AA_TOGGLE</type>
<position>-42,-390.5</position>
<output>
<ID>OUT_0</ID>97 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>260</ID>
<type>AE_OR2</type>
<position>-8.5,-399</position>
<input>
<ID>IN_0</ID>96 </input>
<input>
<ID>IN_1</ID>97 </input>
<output>
<ID>OUT</ID>99 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>262</ID>
<type>AA_AND2</type>
<position>-8,-408.5</position>
<input>
<ID>IN_0</ID>98 </input>
<input>
<ID>IN_1</ID>97 </input>
<output>
<ID>OUT</ID>100 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>264</ID>
<type>GA_LED</type>
<position>-4.5,-399</position>
<input>
<ID>N_in0</ID>99 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>266</ID>
<type>GA_LED</type>
<position>-4,-408.5</position>
<input>
<ID>N_in0</ID>100 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>268</ID>
<type>BA_DECODER_2x4</type>
<position>-48.5,-437</position>
<input>
<ID>ENABLE</ID>101 </input>
<input>
<ID>IN_0</ID>103 </input>
<input>
<ID>IN_1</ID>102 </input>
<output>
<ID>OUT_0</ID>107 </output>
<output>
<ID>OUT_1</ID>106 </output>
<output>
<ID>OUT_2</ID>105 </output>
<output>
<ID>OUT_3</ID>104 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>270</ID>
<type>AA_TOGGLE</type>
<position>-60,-432.5</position>
<output>
<ID>OUT_0</ID>101 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>272</ID>
<type>AA_TOGGLE</type>
<position>-60,-437</position>
<output>
<ID>OUT_0</ID>102 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>274</ID>
<type>AA_TOGGLE</type>
<position>-60,-441.5</position>
<output>
<ID>OUT_0</ID>103 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>276</ID>
<type>GA_LED</type>
<position>-41,-432</position>
<input>
<ID>N_in0</ID>104 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>278</ID>
<type>GA_LED</type>
<position>-35.5,-436</position>
<input>
<ID>N_in0</ID>105 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>280</ID>
<type>GA_LED</type>
<position>-29.5,-438</position>
<input>
<ID>N_in0</ID>106 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>282</ID>
<type>GA_LED</type>
<position>-36,-442</position>
<input>
<ID>N_in0</ID>107 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>284</ID>
<type>BE_DECODER_3x8</type>
<position>2,-434.5</position>
<input>
<ID>ENABLE</ID>108 </input>
<input>
<ID>IN_0</ID>111 </input>
<input>
<ID>IN_1</ID>110 </input>
<input>
<ID>IN_2</ID>109 </input>
<output>
<ID>OUT_0</ID>119 </output>
<output>
<ID>OUT_1</ID>118 </output>
<output>
<ID>OUT_2</ID>117 </output>
<output>
<ID>OUT_3</ID>116 </output>
<output>
<ID>OUT_4</ID>115 </output>
<output>
<ID>OUT_5</ID>114 </output>
<output>
<ID>OUT_6</ID>113 </output>
<output>
<ID>OUT_7</ID>112 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>286</ID>
<type>AA_TOGGLE</type>
<position>-11,-425</position>
<output>
<ID>OUT_0</ID>108 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>288</ID>
<type>AA_TOGGLE</type>
<position>-9.5,-434</position>
<output>
<ID>OUT_0</ID>109 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>290</ID>
<type>AA_TOGGLE</type>
<position>-12.5,-437</position>
<output>
<ID>OUT_0</ID>110 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>292</ID>
<type>AA_TOGGLE</type>
<position>-6,-441.5</position>
<output>
<ID>OUT_0</ID>111 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>294</ID>
<type>GA_LED</type>
<position>7.5,-425</position>
<input>
<ID>N_in0</ID>112 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>296</ID>
<type>GA_LED</type>
<position>10,-431.5</position>
<input>
<ID>N_in0</ID>113 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>298</ID>
<type>GA_LED</type>
<position>14.5,-433</position>
<input>
<ID>N_in0</ID>114 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>300</ID>
<type>GA_LED</type>
<position>28,-434.5</position>
<input>
<ID>N_in0</ID>115 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>302</ID>
<type>GA_LED</type>
<position>21.5,-435.5</position>
<input>
<ID>N_in0</ID>116 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>304</ID>
<type>GA_LED</type>
<position>13.5,-436.5</position>
<input>
<ID>N_in0</ID>117 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>306</ID>
<type>GA_LED</type>
<position>10.5,-437.5</position>
<input>
<ID>N_in0</ID>118 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>308</ID>
<type>GA_LED</type>
<position>10,-440.5</position>
<input>
<ID>N_in0</ID>119 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>310</ID>
<type>BI_DECODER_4x16</type>
<position>-39.5,-467</position>
<input>
<ID>ENABLE</ID>120 </input>
<input>
<ID>IN_0</ID>124 </input>
<input>
<ID>IN_1</ID>123 </input>
<input>
<ID>IN_2</ID>122 </input>
<input>
<ID>IN_3</ID>121 </input>
<output>
<ID>OUT_0</ID>131 </output>
<output>
<ID>OUT_1</ID>132 </output>
<output>
<ID>OUT_10</ID>130 </output>
<output>
<ID>OUT_11</ID>129 </output>
<output>
<ID>OUT_12</ID>128 </output>
<output>
<ID>OUT_13</ID>127 </output>
<output>
<ID>OUT_14</ID>126 </output>
<output>
<ID>OUT_15</ID>125 </output>
<output>
<ID>OUT_2</ID>133 </output>
<output>
<ID>OUT_3</ID>140 </output>
<output>
<ID>OUT_4</ID>139 </output>
<output>
<ID>OUT_5</ID>138 </output>
<output>
<ID>OUT_6</ID>137 </output>
<output>
<ID>OUT_7</ID>136 </output>
<output>
<ID>OUT_8</ID>135 </output>
<output>
<ID>OUT_9</ID>134 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>312</ID>
<type>AA_TOGGLE</type>
<position>-51.5,-453</position>
<output>
<ID>OUT_0</ID>120 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>314</ID>
<type>AA_TOGGLE</type>
<position>-50,-462.5</position>
<output>
<ID>OUT_0</ID>121 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>316</ID>
<type>AA_TOGGLE</type>
<position>-58.5,-472.5</position>
<output>
<ID>OUT_0</ID>122 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>318</ID>
<type>AA_TOGGLE</type>
<position>-71.5,-474</position>
<output>
<ID>OUT_0</ID>123 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>320</ID>
<type>AA_TOGGLE</type>
<position>-47.5,-480.5</position>
<output>
<ID>OUT_0</ID>124 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>322</ID>
<type>GA_LED</type>
<position>-28,-448</position>
<input>
<ID>N_in0</ID>125 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>324</ID>
<type>GA_LED</type>
<position>-15.5,-449.5</position>
<input>
<ID>N_in0</ID>126 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>326</ID>
<type>GA_LED</type>
<position>-12,-451</position>
<input>
<ID>N_in0</ID>127 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>328</ID>
<type>GA_LED</type>
<position>-7,-452.5</position>
<input>
<ID>N_in0</ID>128 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>330</ID>
<type>GA_LED</type>
<position>-2,-454.5</position>
<input>
<ID>N_in0</ID>129 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>332</ID>
<type>GA_LED</type>
<position>-11.5,-456.5</position>
<input>
<ID>N_in0</ID>130 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>334</ID>
<type>GA_LED</type>
<position>-33.5,-483</position>
<input>
<ID>N_in0</ID>131 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>336</ID>
<type>GA_LED</type>
<position>-13,-473.5</position>
<input>
<ID>N_in0</ID>132 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>338</ID>
<type>GA_LED</type>
<position>-9.5,-472</position>
<input>
<ID>N_in0</ID>133 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>340</ID>
<type>GA_LED</type>
<position>-7.5,-459</position>
<input>
<ID>N_in0</ID>134 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>342</ID>
<type>GA_LED</type>
<position>1,-460</position>
<input>
<ID>N_in0</ID>135 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>344</ID>
<type>GA_LED</type>
<position>2,-462.5</position>
<input>
<ID>N_in0</ID>136 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>346</ID>
<type>GA_LED</type>
<position>5,-465</position>
<input>
<ID>N_in0</ID>137 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>348</ID>
<type>GA_LED</type>
<position>9.5,-467</position>
<input>
<ID>N_in0</ID>138 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>350</ID>
<type>GA_LED</type>
<position>16.5,-468.5</position>
<input>
<ID>N_in0</ID>139 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>352</ID>
<type>GA_LED</type>
<position>-25,-470</position>
<input>
<ID>N_in0</ID>140 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>354</ID>
<type>AA_TOGGLE</type>
<position>-56,-495.5</position>
<output>
<ID>OUT_0</ID>143 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>356</ID>
<type>AA_TOGGLE</type>
<position>-56,-502</position>
<output>
<ID>OUT_0</ID>144 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>358</ID>
<type>AA_TOGGLE</type>
<position>-56,-508.5</position>
<output>
<ID>OUT_0</ID>145 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>360</ID>
<type>AA_TOGGLE</type>
<position>-56,-515</position>
<output>
<ID>OUT_0</ID>146 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>362</ID>
<type>AI_XOR2</type>
<position>-41.5,-498</position>
<input>
<ID>IN_0</ID>143 </input>
<input>
<ID>IN_1</ID>144 </input>
<output>
<ID>OUT</ID>149 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>364</ID>
<type>AI_XOR2</type>
<position>-41.5,-505.5</position>
<input>
<ID>IN_0</ID>144 </input>
<input>
<ID>IN_1</ID>145 </input>
<output>
<ID>OUT</ID>148 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>366</ID>
<type>AI_XOR2</type>
<position>-41.5,-512.5</position>
<input>
<ID>IN_0</ID>145 </input>
<input>
<ID>IN_1</ID>146 </input>
<output>
<ID>OUT</ID>147 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>368</ID>
<type>GA_LED</type>
<position>-20.5,-490.5</position>
<input>
<ID>N_in0</ID>143 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>370</ID>
<type>GA_LED</type>
<position>-21,-498</position>
<input>
<ID>N_in0</ID>149 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>372</ID>
<type>GA_LED</type>
<position>-20.5,-504.5</position>
<input>
<ID>N_in0</ID>148 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>374</ID>
<type>GA_LED</type>
<position>-20,-512</position>
<input>
<ID>N_in0</ID>147 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>376</ID>
<type>AA_TOGGLE</type>
<position>-45.5,-528</position>
<output>
<ID>OUT_0</ID>150 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>378</ID>
<type>AA_TOGGLE</type>
<position>-45.5,-535</position>
<output>
<ID>OUT_0</ID>151 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>380</ID>
<type>AA_TOGGLE</type>
<position>-45.5,-542.5</position>
<output>
<ID>OUT_0</ID>156 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>382</ID>
<type>AA_TOGGLE</type>
<position>-45.5,-550</position>
<output>
<ID>OUT_0</ID>153 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>384</ID>
<type>AI_XOR2</type>
<position>-32.5,-532</position>
<input>
<ID>IN_0</ID>150 </input>
<input>
<ID>IN_1</ID>151 </input>
<output>
<ID>OUT</ID>152 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>386</ID>
<type>GA_LED</type>
<position>-9,-526</position>
<input>
<ID>N_in0</ID>150 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>388</ID>
<type>GA_LED</type>
<position>-9,-532.5</position>
<input>
<ID>N_in0</ID>152 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>2</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>18,-10.5,32.5,-10.5</points>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection>
<intersection>32.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>32.5,-11.5,32.5,-10.5</points>
<connection>
<GID>2</GID>
<name>IN_1</name></connection>
<intersection>-10.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32.5,-17,32.5,-13.5</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<intersection>-17 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>18,-17,32.5,-17</points>
<connection>
<GID>8</GID>
<name>OUT_0</name></connection>
<intersection>32.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34.5,-10,34.5,-7</points>
<connection>
<GID>2</GID>
<name>SEL_0</name></connection>
<connection>
<GID>10</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36.5,-12.5,36.5,-12.5</points>
<connection>
<GID>2</GID>
<name>OUT</name></connection>
<connection>
<GID>12</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80,-11.5,80,-9.5</points>
<connection>
<GID>14</GID>
<name>IN_3</name></connection>
<intersection>-9.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>69,-9.5,80,-9.5</points>
<connection>
<GID>16</GID>
<name>OUT_0</name></connection>
<intersection>80 0</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>69,-13.5,80,-13.5</points>
<connection>
<GID>18</GID>
<name>OUT_0</name></connection>
<intersection>80 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>80,-13.5,80,-13.5</points>
<connection>
<GID>14</GID>
<name>IN_2</name></connection>
<intersection>-13.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80,-16,80,-15.5</points>
<connection>
<GID>14</GID>
<name>IN_1</name></connection>
<intersection>-16 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>63,-16,80,-16</points>
<connection>
<GID>20</GID>
<name>OUT_0</name></connection>
<intersection>80 0</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80,-19.5,80,-17.5</points>
<connection>
<GID>14</GID>
<name>IN_0</name></connection>
<intersection>-19.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>69,-19.5,80,-19.5</points>
<connection>
<GID>22</GID>
<name>OUT_0</name></connection>
<intersection>80 0</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>83,-9.5,83,-6.5</points>
<connection>
<GID>14</GID>
<name>SEL_1</name></connection>
<connection>
<GID>24</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90,-9.5,90,-5.5</points>
<connection>
<GID>26</GID>
<name>OUT_0</name></connection>
<intersection>-9.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>84,-9.5,90,-9.5</points>
<connection>
<GID>14</GID>
<name>SEL_0</name></connection>
<intersection>90 0</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>86,-14.5,99.5,-14.5</points>
<connection>
<GID>14</GID>
<name>OUT</name></connection>
<connection>
<GID>28</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32,-38.5,32,-32.5</points>
<connection>
<GID>30</GID>
<name>IN_7</name></connection>
<intersection>-32.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>25.5,-32.5,32,-32.5</points>
<connection>
<GID>32</GID>
<name>OUT_0</name></connection>
<intersection>32 0</intersection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>25.5,-39.5,32,-39.5</points>
<connection>
<GID>30</GID>
<name>IN_6</name></connection>
<connection>
<GID>34</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32,-40.5,32,-36</points>
<connection>
<GID>30</GID>
<name>IN_5</name></connection>
<intersection>-36 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>25.5,-36,32,-36</points>
<connection>
<GID>36</GID>
<name>OUT_0</name></connection>
<intersection>32 0</intersection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32,-42.5,32,-41.5</points>
<connection>
<GID>30</GID>
<name>IN_4</name></connection>
<intersection>-42.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>25,-42.5,32,-42.5</points>
<connection>
<GID>38</GID>
<name>OUT_0</name></connection>
<intersection>32 0</intersection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32,-44,32,-43.5</points>
<connection>
<GID>30</GID>
<name>IN_2</name></connection>
<intersection>-44 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>19,-44,32,-44</points>
<connection>
<GID>40</GID>
<name>OUT_0</name></connection>
<intersection>32 0</intersection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32,-47.5,32,-44.5</points>
<connection>
<GID>30</GID>
<name>IN_1</name></connection>
<intersection>-47.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>23.5,-47.5,32,-47.5</points>
<connection>
<GID>42</GID>
<name>OUT_0</name></connection>
<intersection>32 0</intersection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32,-50,32,-45.5</points>
<connection>
<GID>30</GID>
<name>IN_0</name></connection>
<intersection>-50 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>29.5,-50,32,-50</points>
<connection>
<GID>44</GID>
<name>OUT_0</name></connection>
<intersection>32 0</intersection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32.5,-36.5,32.5,-30.5</points>
<connection>
<GID>46</GID>
<name>OUT_0</name></connection>
<intersection>-36.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>32.5,-36.5,34,-36.5</points>
<connection>
<GID>30</GID>
<name>SEL_2</name></connection>
<intersection>32.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35,-36.5,35,-30.5</points>
<connection>
<GID>30</GID>
<name>SEL_1</name></connection>
<connection>
<GID>48</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38.5,-36.5,38.5,-30.5</points>
<connection>
<GID>50</GID>
<name>OUT_0</name></connection>
<intersection>-36.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>36,-36.5,38.5,-36.5</points>
<connection>
<GID>30</GID>
<name>SEL_0</name></connection>
<intersection>38.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38,-42,38,-42</points>
<connection>
<GID>52</GID>
<name>N_in0</name></connection>
<connection>
<GID>30</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9.5,-63.5,9.5,-62.5</points>
<connection>
<GID>74</GID>
<name>IN_1</name></connection>
<intersection>-62.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>3.5,-62.5,9.5,-62.5</points>
<connection>
<GID>82</GID>
<name>OUT_0</name></connection>
<intersection>9.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>4,-66,9.5,-66</points>
<connection>
<GID>84</GID>
<name>OUT_0</name></connection>
<intersection>9.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>9.5,-66,9.5,-65.5</points>
<connection>
<GID>74</GID>
<name>IN_0</name></connection>
<intersection>-66 1</intersection></vsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9.5,-72,9.5,-71</points>
<connection>
<GID>76</GID>
<name>IN_1</name></connection>
<intersection>-71 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>4,-71,9.5,-71</points>
<connection>
<GID>86</GID>
<name>OUT_0</name></connection>
<intersection>9.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>4,-74.5,9.5,-74.5</points>
<connection>
<GID>88</GID>
<name>OUT_0</name></connection>
<intersection>9.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>9.5,-74.5,9.5,-74</points>
<connection>
<GID>76</GID>
<name>IN_0</name></connection>
<intersection>-74.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9.5,-80.5,9.5,-80</points>
<connection>
<GID>78</GID>
<name>IN_1</name></connection>
<intersection>-80 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>4.5,-80,9.5,-80</points>
<connection>
<GID>90</GID>
<name>OUT_0</name></connection>
<intersection>9.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>4.5,-82.5,9.5,-82.5</points>
<connection>
<GID>78</GID>
<name>IN_0</name></connection>
<connection>
<GID>92</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9.5,-90,9.5,-89</points>
<connection>
<GID>80</GID>
<name>IN_1</name></connection>
<intersection>-89 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>5,-89,9.5,-89</points>
<connection>
<GID>94</GID>
<name>OUT_0</name></connection>
<intersection>9.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9.5,-92.5,9.5,-92</points>
<connection>
<GID>80</GID>
<name>IN_0</name></connection>
<intersection>-92.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>5,-92.5,9.5,-92.5</points>
<connection>
<GID>96</GID>
<name>OUT_0</name></connection>
<intersection>9.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>13.5,-88.5,13.5,-58.5</points>
<connection>
<GID>98</GID>
<name>OUT_0</name></connection>
<intersection>-88.5 1</intersection>
<intersection>-79 4</intersection>
<intersection>-70.5 3</intersection>
<intersection>-62 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>11.5,-88.5,13.5,-88.5</points>
<connection>
<GID>80</GID>
<name>SEL_0</name></connection>
<intersection>13.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>11.5,-62,13.5,-62</points>
<connection>
<GID>74</GID>
<name>SEL_0</name></connection>
<intersection>13.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>11.5,-70.5,13.5,-70.5</points>
<connection>
<GID>76</GID>
<name>SEL_0</name></connection>
<intersection>13.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>11.5,-79,13.5,-79</points>
<connection>
<GID>78</GID>
<name>SEL_0</name></connection>
<intersection>13.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>43.5,-75.5,43.5,-59.5</points>
<connection>
<GID>112</GID>
<name>OUT_0</name></connection>
<intersection>-75.5 1</intersection>
<intersection>-63 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>43,-75.5,43.5,-75.5</points>
<intersection>43 2</intersection>
<intersection>43.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>43,-76,43,-75.5</points>
<connection>
<GID>102</GID>
<name>SEL_0</name></connection>
<intersection>-75.5 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>41.5,-63,43.5,-63</points>
<connection>
<GID>100</GID>
<name>SEL_0</name></connection>
<intersection>43.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>59.5,-69.5,59.5,-59.5</points>
<connection>
<GID>118</GID>
<name>OUT_0</name></connection>
<intersection>-69.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>59.5,-69.5,59.5,-69.5</points>
<connection>
<GID>116</GID>
<name>SEL_0</name></connection>
<intersection>59.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>13.5,-64.5,39.5,-64.5</points>
<connection>
<GID>100</GID>
<name>IN_1</name></connection>
<connection>
<GID>74</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26.5,-73,26.5,-66.5</points>
<intersection>-73 2</intersection>
<intersection>-66.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26.5,-66.5,39.5,-66.5</points>
<connection>
<GID>100</GID>
<name>IN_0</name></connection>
<intersection>26.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>13.5,-73,26.5,-73</points>
<connection>
<GID>76</GID>
<name>OUT</name></connection>
<intersection>26.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26.5,-81.5,26.5,-77.5</points>
<intersection>-81.5 2</intersection>
<intersection>-77.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26.5,-77.5,41,-77.5</points>
<connection>
<GID>102</GID>
<name>IN_1</name></connection>
<intersection>26.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>13.5,-81.5,26.5,-81.5</points>
<connection>
<GID>78</GID>
<name>OUT</name></connection>
<intersection>26.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28.5,-91,28.5,-79.5</points>
<intersection>-91 2</intersection>
<intersection>-79.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>28.5,-79.5,41,-79.5</points>
<connection>
<GID>102</GID>
<name>IN_0</name></connection>
<intersection>28.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>13.5,-91,28.5,-91</points>
<connection>
<GID>80</GID>
<name>OUT</name></connection>
<intersection>28.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>51,-78.5,51,-73</points>
<intersection>-78.5 2</intersection>
<intersection>-73 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>51,-73,57.5,-73</points>
<connection>
<GID>116</GID>
<name>IN_0</name></connection>
<intersection>51 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>45,-78.5,51,-78.5</points>
<connection>
<GID>102</GID>
<name>OUT</name></connection>
<intersection>51 0</intersection></hsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50.5,-71,50.5,-65.5</points>
<intersection>-71 1</intersection>
<intersection>-65.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50.5,-71,57.5,-71</points>
<connection>
<GID>116</GID>
<name>IN_1</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>43.5,-65.5,50.5,-65.5</points>
<connection>
<GID>100</GID>
<name>OUT</name></connection>
<intersection>50.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>46</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>61.5,-72,61.5,-72</points>
<connection>
<GID>120</GID>
<name>N_in0</name></connection>
<connection>
<GID>116</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>48</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>5,-143,5,-101.5</points>
<connection>
<GID>132</GID>
<name>OUT_0</name></connection>
<intersection>-143 3</intersection>
<intersection>-104 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>5,-104,8,-104</points>
<connection>
<GID>138</GID>
<name>IN_0</name></connection>
<intersection>5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>5,-143,41.5,-143</points>
<connection>
<GID>154</GID>
<name>IN_1</name></connection>
<intersection>5 0</intersection>
<intersection>27.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>27.5,-143,27.5,-120</points>
<intersection>-143 3</intersection>
<intersection>-120 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>27.5,-120,41,-120</points>
<connection>
<GID>150</GID>
<name>IN_1</name></connection>
<intersection>27.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>50</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>15,-122,15,-105</points>
<intersection>-122 4</intersection>
<intersection>-109 1</intersection>
<intersection>-105 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>15,-109,40,-109</points>
<connection>
<GID>148</GID>
<name>IN_2</name></connection>
<intersection>15 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-10,-105,15,-105</points>
<connection>
<GID>136</GID>
<name>OUT_0</name></connection>
<intersection>15 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>15,-122,41,-122</points>
<connection>
<GID>150</GID>
<name>IN_2</name></connection>
<intersection>15 0</intersection></hsegment></shape></wire>
<wire>
<ID>52</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>23.5,-105,23.5,-102.5</points>
<connection>
<GID>134</GID>
<name>OUT_0</name></connection>
<intersection>-105 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>23.5,-105,40,-105</points>
<connection>
<GID>148</GID>
<name>IN_0</name></connection>
<intersection>23.5 0</intersection>
<intersection>37.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>37.5,-118,37.5,-105</points>
<intersection>-118 3</intersection>
<intersection>-105 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>37.5,-118,41,-118</points>
<connection>
<GID>150</GID>
<name>IN_0</name></connection>
<intersection>37.5 2</intersection>
<intersection>38.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>38.5,-141,38.5,-118</points>
<intersection>-141 7</intersection>
<intersection>-129.5 5</intersection>
<intersection>-118 3</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>38.5,-129.5,40.5,-129.5</points>
<connection>
<GID>152</GID>
<name>IN_0</name></connection>
<intersection>38.5 4</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>38.5,-141,41.5,-141</points>
<connection>
<GID>154</GID>
<name>IN_0</name></connection>
<intersection>38.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>53</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>46,-107,46,-107</points>
<connection>
<GID>159</GID>
<name>N_in0</name></connection>
<connection>
<GID>148</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>54</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47,-120,47,-120</points>
<connection>
<GID>150</GID>
<name>OUT</name></connection>
<connection>
<GID>161</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>55</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>46.5,-131.5,46.5,-131.5</points>
<connection>
<GID>152</GID>
<name>OUT</name></connection>
<connection>
<GID>163</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>56</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47.5,-143,47.5,-143</points>
<connection>
<GID>154</GID>
<name>OUT</name></connection>
<connection>
<GID>165</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>57</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-16,-145,-16,-101.5</points>
<connection>
<GID>130</GID>
<name>OUT_0</name></connection>
<intersection>-145 5</intersection>
<intersection>-133.5 3</intersection>
<intersection>-105 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-16,-105,-14,-105</points>
<connection>
<GID>136</GID>
<name>IN_0</name></connection>
<intersection>-16 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-16,-133.5,40.5,-133.5</points>
<connection>
<GID>152</GID>
<name>IN_2</name></connection>
<intersection>-16 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-16,-145,41.5,-145</points>
<connection>
<GID>154</GID>
<name>IN_2</name></connection>
<intersection>-16 0</intersection></hsegment></shape></wire>
<wire>
<ID>58</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>21,-131.5,21,-104</points>
<intersection>-131.5 2</intersection>
<intersection>-104 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>12,-104,21,-104</points>
<connection>
<GID>138</GID>
<name>OUT_0</name></connection>
<intersection>21 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>21,-131.5,40.5,-131.5</points>
<connection>
<GID>152</GID>
<name>IN_1</name></connection>
<intersection>21 0</intersection></hsegment></shape></wire>
<wire>
<ID>68</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-11.5,-259,-11.5,-169.5</points>
<connection>
<GID>173</GID>
<name>OUT_0</name></connection>
<intersection>-259 15</intersection>
<intersection>-247 13</intersection>
<intersection>-234.5 11</intersection>
<intersection>-220.5 9</intersection>
<intersection>-205.5 7</intersection>
<intersection>-193.5 5</intersection>
<intersection>-182 3</intersection>
<intersection>-170.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-11.5,-170.5,28,-170.5</points>
<connection>
<GID>175</GID>
<name>IN_0</name></connection>
<intersection>-11.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-11.5,-182,38.5,-182</points>
<connection>
<GID>177</GID>
<name>IN_0</name></connection>
<intersection>-11.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-11.5,-193.5,45.5,-193.5</points>
<connection>
<GID>179</GID>
<name>IN_0</name></connection>
<intersection>-11.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-11.5,-205.5,48,-205.5</points>
<connection>
<GID>181</GID>
<name>IN_0</name></connection>
<intersection>-11.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-11.5,-220.5,39,-220.5</points>
<connection>
<GID>183</GID>
<name>IN_0</name></connection>
<intersection>-11.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>-11.5,-234.5,44,-234.5</points>
<connection>
<GID>185</GID>
<name>IN_0</name></connection>
<intersection>-11.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>-11.5,-247,43,-247</points>
<connection>
<GID>187</GID>
<name>IN_0</name></connection>
<intersection>-11.5 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>-11.5,-259,45.5,-259</points>
<connection>
<GID>189</GID>
<name>IN_0</name></connection>
<intersection>-11.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>69</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-82,-172,-65.5,-172</points>
<connection>
<GID>207</GID>
<name>IN_0</name></connection>
<intersection>-82 5</intersection>
<intersection>-69 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-69,-172,-69,-170</points>
<connection>
<GID>167</GID>
<name>OUT_0</name></connection>
<intersection>-172 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>-82,-238.5,-82,-172</points>
<intersection>-238.5 6</intersection>
<intersection>-226.5 13</intersection>
<intersection>-172 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-82,-238.5,44,-238.5</points>
<connection>
<GID>185</GID>
<name>IN_2</name></connection>
<intersection>-82 5</intersection>
<intersection>-32.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>-32.5,-261,-32.5,-238.5</points>
<intersection>-261 10</intersection>
<intersection>-253 11</intersection>
<intersection>-240.5 12</intersection>
<intersection>-238.5 6</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>-32.5,-261,45.5,-261</points>
<connection>
<GID>189</GID>
<name>IN_1</name></connection>
<intersection>-32.5 7</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>-32.5,-253,43,-253</points>
<connection>
<GID>187</GID>
<name>IN_3</name></connection>
<intersection>-32.5 7</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>-32.5,-240.5,44,-240.5</points>
<connection>
<GID>185</GID>
<name>IN_3</name></connection>
<intersection>-32.5 7</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>-82,-226.5,39,-226.5</points>
<connection>
<GID>183</GID>
<name>IN_3</name></connection>
<intersection>-82 5</intersection></hsegment></shape></wire>
<wire>
<ID>70</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-52,-171,-52,-169.5</points>
<connection>
<GID>169</GID>
<name>OUT_0</name></connection>
<intersection>-171 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-52,-171,-11.5,-171</points>
<connection>
<GID>209</GID>
<name>IN_0</name></connection>
<intersection>-52 0</intersection>
<intersection>-11.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-11.5,-197.5,-11.5,-171</points>
<intersection>-197.5 3</intersection>
<intersection>-171 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-11.5,-197.5,45.5,-197.5</points>
<connection>
<GID>179</GID>
<name>IN_2</name></connection>
<intersection>-11.5 2</intersection>
<intersection>10.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>10.5,-207.5,10.5,-197.5</points>
<intersection>-207.5 5</intersection>
<intersection>-197.5 3</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>10.5,-207.5,48,-207.5</points>
<connection>
<GID>181</GID>
<name>IN_1</name></connection>
<intersection>10.5 4</intersection>
<intersection>15 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>15,-251,15,-207.5</points>
<intersection>-251 7</intersection>
<intersection>-224.5 10</intersection>
<intersection>-207.5 5</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>2,-251,43,-251</points>
<connection>
<GID>187</GID>
<name>IN_2</name></connection>
<intersection>2 8</intersection>
<intersection>15 6</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>2,-263,2,-251</points>
<intersection>-263 9</intersection>
<intersection>-251 7</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>2,-263,45.5,-263</points>
<connection>
<GID>189</GID>
<name>IN_2</name></connection>
<intersection>2 8</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>15,-224.5,39,-224.5</points>
<connection>
<GID>183</GID>
<name>IN_2</name></connection>
<intersection>15 6</intersection></hsegment></shape></wire>
<wire>
<ID>71</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-32.5,-184,-32.5,-169.5</points>
<connection>
<GID>171</GID>
<name>OUT_0</name></connection>
<intersection>-184 3</intersection>
<intersection>-170.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-32.5,-170.5,-30,-170.5</points>
<connection>
<GID>211</GID>
<name>IN_0</name></connection>
<intersection>-32.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-32.5,-184,38.5,-184</points>
<connection>
<GID>177</GID>
<name>IN_1</name></connection>
<intersection>-32.5 0</intersection>
<intersection>6 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>6,-209.5,6,-184</points>
<intersection>-209.5 5</intersection>
<intersection>-184 3</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-57,-209.5,48,-209.5</points>
<connection>
<GID>181</GID>
<name>IN_2</name></connection>
<intersection>-57 6</intersection>
<intersection>6 4</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-57,-265,-57,-209.5</points>
<intersection>-265 8</intersection>
<intersection>-236.5 9</intersection>
<intersection>-209.5 5</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>-57,-265,45.5,-265</points>
<connection>
<GID>189</GID>
<name>IN_3</name></connection>
<intersection>-57 6</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-57,-236.5,44,-236.5</points>
<connection>
<GID>185</GID>
<name>IN_1</name></connection>
<intersection>-57 6</intersection></hsegment></shape></wire>
<wire>
<ID>72</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-6,-172.5,-6,-170.5</points>
<intersection>-172.5 1</intersection>
<intersection>-170.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-17,-172.5,28,-172.5</points>
<connection>
<GID>175</GID>
<name>IN_1</name></connection>
<intersection>-17 3</intersection>
<intersection>-6 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-26,-170.5,-6,-170.5</points>
<connection>
<GID>211</GID>
<name>OUT_0</name></connection>
<intersection>-6 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-17,-195.5,-17,-172.5</points>
<intersection>-195.5 4</intersection>
<intersection>-172.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-44.5,-195.5,45.5,-195.5</points>
<connection>
<GID>179</GID>
<name>IN_1</name></connection>
<intersection>-44.5 5</intersection>
<intersection>-17 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-44.5,-249,-44.5,-195.5</points>
<intersection>-249 6</intersection>
<intersection>-222.5 7</intersection>
<intersection>-195.5 4</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-44.5,-249,43,-249</points>
<connection>
<GID>187</GID>
<name>IN_1</name></connection>
<intersection>-44.5 5</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-44.5,-222.5,39,-222.5</points>
<connection>
<GID>183</GID>
<name>IN_1</name></connection>
<intersection>-44.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>73</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-15,-174.5,-15,-171</points>
<intersection>-174.5 1</intersection>
<intersection>-171 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-15,-174.5,28,-174.5</points>
<connection>
<GID>175</GID>
<name>IN_2</name></connection>
<intersection>-15 0</intersection>
<intersection>8 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-44.5,-171,-15,-171</points>
<connection>
<GID>209</GID>
<name>OUT_0</name></connection>
<intersection>-15 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>8,-186,8,-174.5</points>
<intersection>-186 4</intersection>
<intersection>-174.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>8,-186,38.5,-186</points>
<connection>
<GID>177</GID>
<name>IN_2</name></connection>
<intersection>8 3</intersection></hsegment></shape></wire>
<wire>
<ID>74</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-23.5,-176.5,-23.5,-172</points>
<intersection>-176.5 1</intersection>
<intersection>-172 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-28,-176.5,28,-176.5</points>
<connection>
<GID>175</GID>
<name>IN_3</name></connection>
<intersection>-28 3</intersection>
<intersection>-23.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-61.5,-172,-23.5,-172</points>
<connection>
<GID>207</GID>
<name>OUT_0</name></connection>
<intersection>-23.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-28,-199.5,-28,-176.5</points>
<intersection>-199.5 6</intersection>
<intersection>-188 4</intersection>
<intersection>-176.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-28,-188,38.5,-188</points>
<connection>
<GID>177</GID>
<name>IN_3</name></connection>
<intersection>-28 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-28,-199.5,45.5,-199.5</points>
<connection>
<GID>179</GID>
<name>IN_3</name></connection>
<intersection>-28 3</intersection>
<intersection>-11.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>-11.5,-211.5,-11.5,-199.5</points>
<intersection>-211.5 8</intersection>
<intersection>-199.5 6</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>-11.5,-211.5,48,-211.5</points>
<connection>
<GID>181</GID>
<name>IN_3</name></connection>
<intersection>-11.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>75</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>51.5,-262,51.5,-262</points>
<connection>
<GID>212</GID>
<name>N_in0</name></connection>
<connection>
<GID>189</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>76</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49,-250,49,-250</points>
<connection>
<GID>213</GID>
<name>N_in0</name></connection>
<connection>
<GID>187</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>77</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50,-237.5,50,-237.5</points>
<connection>
<GID>214</GID>
<name>N_in0</name></connection>
<connection>
<GID>185</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>78</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>45,-223.5,45,-223.5</points>
<connection>
<GID>215</GID>
<name>N_in0</name></connection>
<connection>
<GID>183</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>79</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54,-208.5,54,-208.5</points>
<connection>
<GID>181</GID>
<name>OUT</name></connection>
<connection>
<GID>216</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>80</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>51.5,-196.5,51.5,-196.5</points>
<connection>
<GID>179</GID>
<name>OUT</name></connection>
<connection>
<GID>218</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>81</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>44.5,-185,44.5,-185</points>
<connection>
<GID>177</GID>
<name>OUT</name></connection>
<connection>
<GID>219</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>82</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34,-173.5,34,-173.5</points>
<connection>
<GID>175</GID>
<name>OUT</name></connection>
<connection>
<GID>220</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>83</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-10.5,-304,-10.5,-299.5</points>
<connection>
<GID>236</GID>
<name>OUT_0</name></connection>
<intersection>-304 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-11,-304,29.5,-304</points>
<connection>
<GID>238</GID>
<name>IN_0</name></connection>
<intersection>-11 2</intersection>
<intersection>-10.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-11,-340,-11,-304</points>
<intersection>-340 3</intersection>
<intersection>-304 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-11,-340,30,-340</points>
<connection>
<GID>242</GID>
<name>IN_3</name></connection>
<intersection>-11 2</intersection>
<intersection>14 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>14,-367.5,14,-340</points>
<intersection>-367.5 5</intersection>
<intersection>-340 3</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>14,-367.5,31,-367.5</points>
<connection>
<GID>244</GID>
<name>IN_3</name></connection>
<intersection>14 4</intersection></hsegment></shape></wire>
<wire>
<ID>84</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-23.5,-306,-23.5,-299</points>
<connection>
<GID>234</GID>
<name>OUT_0</name></connection>
<intersection>-306 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-23.5,-306,29.5,-306</points>
<connection>
<GID>238</GID>
<name>IN_1</name></connection>
<intersection>-23.5 0</intersection>
<intersection>14 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>14,-338,14,-306</points>
<intersection>-338 3</intersection>
<intersection>-306 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>14,-338,30,-338</points>
<connection>
<GID>242</GID>
<name>IN_2</name></connection>
<intersection>14 2</intersection></hsegment></shape></wire>
<wire>
<ID>85</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-33,-365.5,-33,-299</points>
<connection>
<GID>232</GID>
<name>OUT_0</name></connection>
<intersection>-365.5 3</intersection>
<intersection>-308 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-33,-308,29.5,-308</points>
<connection>
<GID>238</GID>
<name>IN_2</name></connection>
<intersection>-33 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-33,-365.5,31,-365.5</points>
<connection>
<GID>244</GID>
<name>IN_2</name></connection>
<intersection>-33 0</intersection></hsegment></shape></wire>
<wire>
<ID>86</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-43.5,-310,-43.5,-299.5</points>
<connection>
<GID>230</GID>
<name>OUT_0</name></connection>
<intersection>-310 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-43.5,-310,29.5,-310</points>
<connection>
<GID>238</GID>
<name>IN_3</name></connection>
<intersection>-43.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>87</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-64.5,-334,-64.5,-299</points>
<connection>
<GID>226</GID>
<name>OUT_0</name></connection>
<intersection>-334 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-64.5,-334,30,-334</points>
<connection>
<GID>242</GID>
<name>IN_0</name></connection>
<intersection>-64.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>88</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-54.5,-336,-54.5,-299.5</points>
<connection>
<GID>228</GID>
<name>OUT_0</name></connection>
<intersection>-336 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-54.5,-336,30,-336</points>
<connection>
<GID>242</GID>
<name>IN_1</name></connection>
<intersection>-54.5 0</intersection>
<intersection>6 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>6,-363.5,6,-336</points>
<intersection>-363.5 3</intersection>
<intersection>-336 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>6,-363.5,31,-363.5</points>
<connection>
<GID>244</GID>
<name>IN_1</name></connection>
<intersection>6 2</intersection></hsegment></shape></wire>
<wire>
<ID>90</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-77.5,-361.5,-77.5,-299.5</points>
<connection>
<GID>224</GID>
<name>OUT_0</name></connection>
<intersection>-361.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-77.5,-361.5,31,-361.5</points>
<connection>
<GID>244</GID>
<name>IN_0</name></connection>
<intersection>-77.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>91</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36.5,-307,36.5,-307</points>
<connection>
<GID>238</GID>
<name>OUT</name></connection>
<connection>
<GID>246</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>92</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37,-337,37,-337</points>
<connection>
<GID>242</GID>
<name>OUT</name></connection>
<connection>
<GID>248</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>93</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38,-364.5,38,-364.5</points>
<connection>
<GID>244</GID>
<name>OUT</name></connection>
<connection>
<GID>250</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>96</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-56,-398,-56,-392.5</points>
<connection>
<GID>256</GID>
<name>OUT_0</name></connection>
<intersection>-398 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-56,-398,-11.5,-398</points>
<connection>
<GID>260</GID>
<name>IN_0</name></connection>
<intersection>-56 0</intersection></hsegment></shape></wire>
<wire>
<ID>97</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-42,-400,-42,-392.5</points>
<connection>
<GID>258</GID>
<name>OUT_0</name></connection>
<intersection>-400 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-42,-400,-11.5,-400</points>
<connection>
<GID>260</GID>
<name>IN_1</name></connection>
<intersection>-42 0</intersection>
<intersection>-28 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-28,-410,-28,-400</points>
<intersection>-410 3</intersection>
<intersection>-400 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-28,-410,-11,-410</points>
<intersection>-28 2</intersection>
<intersection>-11 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-11,-410,-11,-409.5</points>
<connection>
<GID>262</GID>
<name>IN_1</name></connection>
<intersection>-410 3</intersection></vsegment></shape></wire>
<wire>
<ID>98</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-70,-407.5,-70,-392.5</points>
<connection>
<GID>254</GID>
<name>OUT_0</name></connection>
<intersection>-407.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-70,-407.5,-11,-407.5</points>
<connection>
<GID>262</GID>
<name>IN_0</name></connection>
<intersection>-70 0</intersection></hsegment></shape></wire>
<wire>
<ID>99</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-5.5,-399,-5.5,-399</points>
<connection>
<GID>260</GID>
<name>OUT</name></connection>
<connection>
<GID>264</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>100</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-5,-408.5,-5,-408.5</points>
<connection>
<GID>262</GID>
<name>OUT</name></connection>
<connection>
<GID>266</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>101</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-51.5,-435.5,-51.5,-432.5</points>
<connection>
<GID>268</GID>
<name>ENABLE</name></connection>
<intersection>-432.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-58,-432.5,-51.5,-432.5</points>
<connection>
<GID>270</GID>
<name>OUT_0</name></connection>
<intersection>-51.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>102</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-51.5,-437.5,-51.5,-437</points>
<connection>
<GID>268</GID>
<name>IN_1</name></connection>
<intersection>-437 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-58,-437,-51.5,-437</points>
<connection>
<GID>272</GID>
<name>OUT_0</name></connection>
<intersection>-51.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>103</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-51.5,-441.5,-51.5,-438.5</points>
<connection>
<GID>268</GID>
<name>IN_0</name></connection>
<intersection>-441.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-58,-441.5,-51.5,-441.5</points>
<connection>
<GID>274</GID>
<name>OUT_0</name></connection>
<intersection>-51.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>104</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-45.5,-435.5,-45.5,-432</points>
<connection>
<GID>268</GID>
<name>OUT_3</name></connection>
<intersection>-432 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-45.5,-432,-42,-432</points>
<connection>
<GID>276</GID>
<name>N_in0</name></connection>
<intersection>-45.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>105</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-45.5,-436,-36.5,-436</points>
<connection>
<GID>278</GID>
<name>N_in0</name></connection>
<intersection>-45.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-45.5,-436.5,-45.5,-436</points>
<connection>
<GID>268</GID>
<name>OUT_2</name></connection>
<intersection>-436 1</intersection></vsegment></shape></wire>
<wire>
<ID>106</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-45.5,-438,-45.5,-437.5</points>
<connection>
<GID>268</GID>
<name>OUT_1</name></connection>
<intersection>-438 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-45.5,-438,-30.5,-438</points>
<connection>
<GID>280</GID>
<name>N_in0</name></connection>
<intersection>-45.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>107</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-45.5,-442,-45.5,-438.5</points>
<connection>
<GID>268</GID>
<name>OUT_0</name></connection>
<intersection>-442 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-45.5,-442,-37,-442</points>
<connection>
<GID>282</GID>
<name>N_in0</name></connection>
<intersection>-45.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>108</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1,-431,-1,-425</points>
<connection>
<GID>284</GID>
<name>ENABLE</name></connection>
<intersection>-425 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-9,-425,-1,-425</points>
<connection>
<GID>286</GID>
<name>OUT_0</name></connection>
<intersection>-1 0</intersection></hsegment></shape></wire>
<wire>
<ID>109</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1,-436,-1,-434</points>
<connection>
<GID>284</GID>
<name>IN_2</name></connection>
<intersection>-434 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-7.5,-434,-1,-434</points>
<connection>
<GID>288</GID>
<name>OUT_0</name></connection>
<intersection>-1 0</intersection></hsegment></shape></wire>
<wire>
<ID>110</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-10.5,-437,-1,-437</points>
<connection>
<GID>284</GID>
<name>IN_1</name></connection>
<connection>
<GID>290</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>111</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1,-441.5,-1,-438</points>
<connection>
<GID>284</GID>
<name>IN_0</name></connection>
<intersection>-441.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-4,-441.5,-1,-441.5</points>
<connection>
<GID>292</GID>
<name>OUT_0</name></connection>
<intersection>-1 0</intersection></hsegment></shape></wire>
<wire>
<ID>112</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>5,-431,5,-425</points>
<connection>
<GID>284</GID>
<name>OUT_7</name></connection>
<intersection>-425 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>5,-425,6.5,-425</points>
<connection>
<GID>294</GID>
<name>N_in0</name></connection>
<intersection>5 0</intersection></hsegment></shape></wire>
<wire>
<ID>113</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>5,-432,5,-431.5</points>
<connection>
<GID>284</GID>
<name>OUT_6</name></connection>
<intersection>-431.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>5,-431.5,9,-431.5</points>
<connection>
<GID>296</GID>
<name>N_in0</name></connection>
<intersection>5 0</intersection></hsegment></shape></wire>
<wire>
<ID>114</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>5,-433,13.5,-433</points>
<connection>
<GID>284</GID>
<name>OUT_5</name></connection>
<connection>
<GID>298</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>115</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>5,-434.5,5,-434</points>
<connection>
<GID>284</GID>
<name>OUT_4</name></connection>
<intersection>-434.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>5,-434.5,27,-434.5</points>
<connection>
<GID>300</GID>
<name>N_in0</name></connection>
<intersection>5 0</intersection></hsegment></shape></wire>
<wire>
<ID>116</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>5,-435.5,20.5,-435.5</points>
<connection>
<GID>302</GID>
<name>N_in0</name></connection>
<intersection>5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>5,-435.5,5,-435</points>
<connection>
<GID>284</GID>
<name>OUT_3</name></connection>
<intersection>-435.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>117</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>5,-436.5,5,-436</points>
<connection>
<GID>284</GID>
<name>OUT_2</name></connection>
<intersection>-436.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>5,-436.5,12.5,-436.5</points>
<connection>
<GID>304</GID>
<name>N_in0</name></connection>
<intersection>5 0</intersection></hsegment></shape></wire>
<wire>
<ID>118</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>5,-437.5,5,-437</points>
<connection>
<GID>284</GID>
<name>OUT_1</name></connection>
<intersection>-437.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>5,-437.5,9.5,-437.5</points>
<connection>
<GID>306</GID>
<name>N_in0</name></connection>
<intersection>5 0</intersection></hsegment></shape></wire>
<wire>
<ID>119</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>5,-440.5,5,-438</points>
<connection>
<GID>284</GID>
<name>OUT_0</name></connection>
<intersection>-440.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>5,-440.5,9,-440.5</points>
<connection>
<GID>308</GID>
<name>N_in0</name></connection>
<intersection>5 0</intersection></hsegment></shape></wire>
<wire>
<ID>120</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-42.5,-459.5,-42.5,-453</points>
<connection>
<GID>310</GID>
<name>ENABLE</name></connection>
<intersection>-453 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-49.5,-453,-42.5,-453</points>
<connection>
<GID>312</GID>
<name>OUT_0</name></connection>
<intersection>-42.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>121</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-42.5,-471.5,-42.5,-462.5</points>
<connection>
<GID>310</GID>
<name>IN_3</name></connection>
<intersection>-462.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-48,-462.5,-42.5,-462.5</points>
<connection>
<GID>314</GID>
<name>OUT_0</name></connection>
<intersection>-42.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>122</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-56.5,-472.5,-42.5,-472.5</points>
<connection>
<GID>310</GID>
<name>IN_2</name></connection>
<connection>
<GID>316</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>123</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-42.5,-474,-42.5,-473.5</points>
<connection>
<GID>310</GID>
<name>IN_1</name></connection>
<intersection>-474 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-69.5,-474,-42.5,-474</points>
<connection>
<GID>318</GID>
<name>OUT_0</name></connection>
<intersection>-42.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>124</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-42.5,-480.5,-42.5,-474.5</points>
<connection>
<GID>310</GID>
<name>IN_0</name></connection>
<intersection>-480.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-45.5,-480.5,-42.5,-480.5</points>
<connection>
<GID>320</GID>
<name>OUT_0</name></connection>
<intersection>-42.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>125</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-36.5,-459.5,-36.5,-448</points>
<connection>
<GID>310</GID>
<name>OUT_15</name></connection>
<intersection>-448 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-36.5,-448,-29,-448</points>
<connection>
<GID>322</GID>
<name>N_in0</name></connection>
<intersection>-36.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>126</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-36.5,-460.5,-36.5,-449.5</points>
<connection>
<GID>310</GID>
<name>OUT_14</name></connection>
<intersection>-449.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-36.5,-449.5,-16.5,-449.5</points>
<connection>
<GID>324</GID>
<name>N_in0</name></connection>
<intersection>-36.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>127</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-36.5,-461.5,-36.5,-451</points>
<connection>
<GID>310</GID>
<name>OUT_13</name></connection>
<intersection>-451 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-36.5,-451,-13,-451</points>
<connection>
<GID>326</GID>
<name>N_in0</name></connection>
<intersection>-36.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>128</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-36.5,-462.5,-36.5,-452.5</points>
<connection>
<GID>310</GID>
<name>OUT_12</name></connection>
<intersection>-452.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-36.5,-452.5,-8,-452.5</points>
<connection>
<GID>328</GID>
<name>N_in0</name></connection>
<intersection>-36.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>129</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-36.5,-454.5,-3,-454.5</points>
<connection>
<GID>330</GID>
<name>N_in0</name></connection>
<intersection>-36.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-36.5,-463.5,-36.5,-454.5</points>
<connection>
<GID>310</GID>
<name>OUT_11</name></connection>
<intersection>-454.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>130</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-36.5,-464.5,-36.5,-456.5</points>
<connection>
<GID>310</GID>
<name>OUT_10</name></connection>
<intersection>-456.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-36.5,-456.5,-12.5,-456.5</points>
<connection>
<GID>332</GID>
<name>N_in0</name></connection>
<intersection>-36.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>131</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-36.5,-483,-36.5,-474.5</points>
<connection>
<GID>310</GID>
<name>OUT_0</name></connection>
<intersection>-483 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-36.5,-483,-34.5,-483</points>
<connection>
<GID>334</GID>
<name>N_in0</name></connection>
<intersection>-36.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>132</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-36.5,-473.5,-14,-473.5</points>
<connection>
<GID>310</GID>
<name>OUT_1</name></connection>
<connection>
<GID>336</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>133</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-36.5,-472.5,-36.5,-472</points>
<connection>
<GID>310</GID>
<name>OUT_2</name></connection>
<intersection>-472 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-36.5,-472,-10.5,-472</points>
<connection>
<GID>338</GID>
<name>N_in0</name></connection>
<intersection>-36.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>134</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-36.5,-465.5,-36.5,-459</points>
<connection>
<GID>310</GID>
<name>OUT_9</name></connection>
<intersection>-459 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-36.5,-459,-8.5,-459</points>
<connection>
<GID>340</GID>
<name>N_in0</name></connection>
<intersection>-36.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>135</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-36.5,-461.5,-5.5,-461.5</points>
<intersection>-36.5 3</intersection>
<intersection>-5.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-5.5,-461.5,-5.5,-460</points>
<intersection>-461.5 1</intersection>
<intersection>-460 4</intersection></vsegment>
<vsegment>
<ID>3</ID>
<points>-36.5,-466.5,-36.5,-461.5</points>
<connection>
<GID>310</GID>
<name>OUT_8</name></connection>
<intersection>-461.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-5.5,-460,0,-460</points>
<connection>
<GID>342</GID>
<name>N_in0</name></connection>
<intersection>-5.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>136</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-36.5,-462.5,1,-462.5</points>
<connection>
<GID>344</GID>
<name>N_in0</name></connection>
<intersection>-36.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-36.5,-467.5,-36.5,-462.5</points>
<connection>
<GID>310</GID>
<name>OUT_7</name></connection>
<intersection>-462.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>137</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-36.5,-468.5,-36.5,-465</points>
<connection>
<GID>310</GID>
<name>OUT_6</name></connection>
<intersection>-465 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-36.5,-465,4,-465</points>
<connection>
<GID>346</GID>
<name>N_in0</name></connection>
<intersection>-36.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>138</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-36.5,-469.5,-36.5,-467</points>
<connection>
<GID>310</GID>
<name>OUT_5</name></connection>
<intersection>-467 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-36.5,-467,8.5,-467</points>
<connection>
<GID>348</GID>
<name>N_in0</name></connection>
<intersection>-36.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>139</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-36.5,-470.5,-36.5,-468.5</points>
<connection>
<GID>310</GID>
<name>OUT_4</name></connection>
<intersection>-468.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-36.5,-468.5,15.5,-468.5</points>
<connection>
<GID>350</GID>
<name>N_in0</name></connection>
<intersection>-36.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>140</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-36.5,-471.5,-36.5,-470</points>
<connection>
<GID>310</GID>
<name>OUT_3</name></connection>
<intersection>-470 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-36.5,-470,-26,-470</points>
<connection>
<GID>352</GID>
<name>N_in0</name></connection>
<intersection>-36.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>143</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-37.5,-495.5,-37.5,-490.5</points>
<intersection>-495.5 2</intersection>
<intersection>-490.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-37.5,-490.5,-21.5,-490.5</points>
<connection>
<GID>368</GID>
<name>N_in0</name></connection>
<intersection>-37.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-54,-495.5,-37.5,-495.5</points>
<connection>
<GID>354</GID>
<name>OUT_0</name></connection>
<intersection>-44.5 3</intersection>
<intersection>-37.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-44.5,-497,-44.5,-495.5</points>
<connection>
<GID>362</GID>
<name>IN_0</name></connection>
<intersection>-495.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>144</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-49,-504.5,-49,-499</points>
<intersection>-504.5 3</intersection>
<intersection>-502 1</intersection>
<intersection>-499 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-54,-502,-49,-502</points>
<connection>
<GID>356</GID>
<name>OUT_0</name></connection>
<intersection>-49 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-49,-499,-44.5,-499</points>
<connection>
<GID>362</GID>
<name>IN_1</name></connection>
<intersection>-49 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-49,-504.5,-44.5,-504.5</points>
<connection>
<GID>364</GID>
<name>IN_0</name></connection>
<intersection>-49 0</intersection></hsegment></shape></wire>
<wire>
<ID>145</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-49,-508.5,-49,-506.5</points>
<intersection>-508.5 1</intersection>
<intersection>-506.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-54,-508.5,-49,-508.5</points>
<connection>
<GID>358</GID>
<name>OUT_0</name></connection>
<intersection>-49 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-49,-506.5,-44.5,-506.5</points>
<connection>
<GID>364</GID>
<name>IN_1</name></connection>
<intersection>-49 0</intersection>
<intersection>-44.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-44.5,-511.5,-44.5,-506.5</points>
<connection>
<GID>366</GID>
<name>IN_0</name></connection>
<intersection>-506.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>146</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-49,-515,-49,-513.5</points>
<intersection>-515 1</intersection>
<intersection>-513.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-54,-515,-49,-515</points>
<connection>
<GID>360</GID>
<name>OUT_0</name></connection>
<intersection>-49 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-49,-513.5,-44.5,-513.5</points>
<connection>
<GID>366</GID>
<name>IN_1</name></connection>
<intersection>-49 0</intersection></hsegment></shape></wire>
<wire>
<ID>147</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-29.5,-512.5,-29.5,-512</points>
<intersection>-512.5 2</intersection>
<intersection>-512 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-29.5,-512,-21,-512</points>
<connection>
<GID>374</GID>
<name>N_in0</name></connection>
<intersection>-29.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-38.5,-512.5,-29.5,-512.5</points>
<connection>
<GID>366</GID>
<name>OUT</name></connection>
<intersection>-29.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>148</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-30,-505.5,-30,-504.5</points>
<intersection>-505.5 2</intersection>
<intersection>-504.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-30,-504.5,-21.5,-504.5</points>
<connection>
<GID>372</GID>
<name>N_in0</name></connection>
<intersection>-30 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-38.5,-505.5,-30,-505.5</points>
<connection>
<GID>364</GID>
<name>OUT</name></connection>
<intersection>-30 0</intersection></hsegment></shape></wire>
<wire>
<ID>149</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-38.5,-498,-22,-498</points>
<connection>
<GID>370</GID>
<name>N_in0</name></connection>
<connection>
<GID>362</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>150</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-26.5,-528,-26.5,-526</points>
<intersection>-528 2</intersection>
<intersection>-526 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-26.5,-526,-10,-526</points>
<connection>
<GID>386</GID>
<name>N_in0</name></connection>
<intersection>-26.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-43.5,-528,-26.5,-528</points>
<connection>
<GID>376</GID>
<name>OUT_0</name></connection>
<intersection>-35.5 3</intersection>
<intersection>-26.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-35.5,-531,-35.5,-528</points>
<connection>
<GID>384</GID>
<name>IN_0</name></connection>
<intersection>-528 2</intersection></vsegment></shape></wire>
<wire>
<ID>151</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-39.5,-535,-39.5,-533</points>
<intersection>-535 2</intersection>
<intersection>-533 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-39.5,-533,-35.5,-533</points>
<connection>
<GID>384</GID>
<name>IN_1</name></connection>
<intersection>-39.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-43.5,-535,-39.5,-535</points>
<connection>
<GID>378</GID>
<name>OUT_0</name></connection>
<intersection>-39.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>152</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-19.5,-532.5,-19.5,-532</points>
<intersection>-532.5 1</intersection>
<intersection>-532 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-19.5,-532.5,-10,-532.5</points>
<connection>
<GID>388</GID>
<name>N_in0</name></connection>
<intersection>-19.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-29.5,-532,-19.5,-532</points>
<connection>
<GID>384</GID>
<name>OUT</name></connection>
<intersection>-27.5 3</intersection>
<intersection>-19.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-27.5,-539.5,-27.5,-532</points>
<connection>
<GID>394</GID>
<name>IN_0</name></connection>
<intersection>-532 2</intersection></vsegment></shape></wire>
<wire>
<ID>153</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-43.5,-550,-20,-550</points>
<connection>
<GID>396</GID>
<name>IN_1</name></connection>
<connection>
<GID>382</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>154</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-15.5,-541.5,-15.5,-540.5</points>
<intersection>-541.5 1</intersection>
<intersection>-540.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-15.5,-541.5,-10,-541.5</points>
<connection>
<GID>390</GID>
<name>N_in0</name></connection>
<intersection>-15.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-21.5,-540.5,-15.5,-540.5</points>
<connection>
<GID>394</GID>
<name>OUT</name></connection>
<intersection>-20 3</intersection>
<intersection>-15.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-20,-548,-20,-540.5</points>
<connection>
<GID>396</GID>
<name>IN_0</name></connection>
<intersection>-540.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>155</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-14,-549,-10,-549</points>
<connection>
<GID>392</GID>
<name>N_in0</name></connection>
<connection>
<GID>396</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>156</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-35.5,-542.5,-35.5,-541.5</points>
<intersection>-542.5 2</intersection>
<intersection>-541.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-35.5,-541.5,-27.5,-541.5</points>
<connection>
<GID>394</GID>
<name>IN_1</name></connection>
<intersection>-35.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-43.5,-542.5,-35.5,-542.5</points>
<connection>
<GID>380</GID>
<name>OUT_0</name></connection>
<intersection>-35.5 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 1>
<page 2>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 2>
<page 3>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 3>
<page 4>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 4>
<page 5>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 5>
<page 6>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 6>
<page 7>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 7>
<page 8>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 8>
<page 9>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 9></circuit>