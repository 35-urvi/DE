<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>34.2741,-268.394,180.074,-342.094</PageViewport>
<gate>
<ID>389</ID>
<type>BA_NAND2</type>
<position>38.5,-205</position>
<input>
<ID>IN_0</ID>206 </input>
<input>
<ID>IN_1</ID>206 </input>
<output>
<ID>OUT</ID>212 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>390</ID>
<type>BA_NAND2</type>
<position>51,-212</position>
<input>
<ID>IN_0</ID>215 </input>
<input>
<ID>IN_1</ID>212 </input>
<output>
<ID>OUT</ID>207 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>391</ID>
<type>BA_NAND2</type>
<position>51,-217</position>
<input>
<ID>IN_0</ID>211 </input>
<input>
<ID>IN_1</ID>206 </input>
<output>
<ID>OUT</ID>208 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2</ID>
<type>AA_AND2</type>
<position>30.5,-14</position>
<input>
<ID>IN_0</ID>2 </input>
<input>
<ID>IN_1</ID>3 </input>
<output>
<ID>OUT</ID>4 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>392</ID>
<type>BA_NAND2</type>
<position>51.5,-225</position>
<input>
<ID>IN_0</ID>211 </input>
<input>
<ID>IN_1</ID>206 </input>
<output>
<ID>OUT</ID>209 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>393</ID>
<type>BA_NAND2</type>
<position>62.5,-225</position>
<input>
<ID>IN_0</ID>209 </input>
<input>
<ID>IN_1</ID>209 </input>
<output>
<ID>OUT</ID>214 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4</ID>
<type>AA_TOGGLE</type>
<position>23,-13</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>394</ID>
<type>BA_NAND2</type>
<position>62.5,-214.5</position>
<input>
<ID>IN_0</ID>207 </input>
<input>
<ID>IN_1</ID>208 </input>
<output>
<ID>OUT</ID>213 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>395</ID>
<type>GA_LED</type>
<position>69.5,-214.5</position>
<input>
<ID>N_in0</ID>213 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>6</ID>
<type>AA_TOGGLE</type>
<position>23,-15</position>
<output>
<ID>OUT_0</ID>3 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>396</ID>
<type>GA_LED</type>
<position>70,-225</position>
<input>
<ID>N_in0</ID>214 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>8</ID>
<type>GA_LED</type>
<position>37.5,-14</position>
<input>
<ID>N_in0</ID>4 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>399</ID>
<type>AA_LABEL</type>
<position>70.5,-211.5</position>
<gparam>LABEL_TEXT diff=ab'+a'b</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>10</ID>
<type>AE_OR2</type>
<position>30.5,-8.5</position>
<input>
<ID>IN_0</ID>9 </input>
<input>
<ID>IN_1</ID>10 </input>
<output>
<ID>OUT</ID>13 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>400</ID>
<type>AA_LABEL</type>
<position>70.5,-222</position>
<gparam>LABEL_TEXT borrow=a'b</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>401</ID>
<type>AA_TOGGLE</type>
<position>89,-200</position>
<output>
<ID>OUT_0</ID>219 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>12</ID>
<type>AA_LABEL</type>
<position>21,-12.5</position>
<gparam>LABEL_TEXT a</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>402</ID>
<type>AA_LABEL</type>
<position>88.5,-197.5</position>
<gparam>LABEL_TEXT a</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>403</ID>
<type>AA_LABEL</type>
<position>98.5,-197.5</position>
<gparam>LABEL_TEXT b</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>404</ID>
<type>BE_NOR2</type>
<position>116,-211.5</position>
<input>
<ID>IN_0</ID>225 </input>
<input>
<ID>IN_1</ID>217 </input>
<output>
<ID>OUT</ID>220 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>405</ID>
<type>BE_NOR2</type>
<position>116,-216.5</position>
<input>
<ID>IN_0</ID>219 </input>
<input>
<ID>IN_1</ID>218 </input>
<output>
<ID>OUT</ID>221 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>16</ID>
<type>AA_LABEL</type>
<position>21,-15</position>
<gparam>LABEL_TEXT b</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>406</ID>
<type>BE_NOR2</type>
<position>115.5,-225.5</position>
<input>
<ID>IN_0</ID>219 </input>
<input>
<ID>IN_1</ID>218 </input>
<output>
<ID>OUT</ID>222 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>407</ID>
<type>BE_NOR2</type>
<position>126,-214</position>
<input>
<ID>IN_0</ID>220 </input>
<input>
<ID>IN_1</ID>221 </input>
<output>
<ID>OUT</ID>224 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>18</ID>
<type>AA_LABEL</type>
<position>41.5,-13.5</position>
<gparam>LABEL_TEXT y=a.b</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>408</ID>
<type>BE_NOR2</type>
<position>93,-207</position>
<input>
<ID>IN_0</ID>219 </input>
<input>
<ID>IN_1</ID>219 </input>
<output>
<ID>OUT</ID>225 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>409</ID>
<type>AA_TOGGLE</type>
<position>98.5,-200</position>
<output>
<ID>OUT_0</ID>217 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>20</ID>
<type>AA_INVERTER</type>
<position>30.5,-3</position>
<input>
<ID>IN_0</ID>11 </input>
<output>
<ID>OUT_0</ID>12 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>410</ID>
<type>BE_NOR2</type>
<position>102.5,-207</position>
<input>
<ID>IN_0</ID>217 </input>
<input>
<ID>IN_1</ID>217 </input>
<output>
<ID>OUT</ID>218 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>411</ID>
<type>GA_LED</type>
<position>141,-214</position>
<input>
<ID>N_in0</ID>223 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>22</ID>
<type>BA_NAND2</type>
<position>59.5,-14.5</position>
<input>
<ID>IN_0</ID>7 </input>
<input>
<ID>IN_1</ID>8 </input>
<output>
<ID>OUT</ID>16 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>412</ID>
<type>GA_LED</type>
<position>123.5,-225.5</position>
<input>
<ID>N_in0</ID>222 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>24</ID>
<type>BE_NOR2</type>
<position>59.5,-9</position>
<input>
<ID>IN_0</ID>5 </input>
<input>
<ID>IN_1</ID>6 </input>
<output>
<ID>OUT</ID>14 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>414</ID>
<type>BE_NOR2</type>
<position>134.5,-214</position>
<input>
<ID>IN_0</ID>224 </input>
<input>
<ID>IN_1</ID>224 </input>
<output>
<ID>OUT</ID>223 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>25</ID>
<type>AA_TOGGLE</type>
<position>52,-10</position>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>26</ID>
<type>AA_TOGGLE</type>
<position>52,-8</position>
<output>
<ID>OUT_0</ID>5 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>416</ID>
<type>AA_LABEL</type>
<position>141.5,-211</position>
<gparam>LABEL_TEXT diff=ab'+a'b</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>27</ID>
<type>AA_TOGGLE</type>
<position>52,-13.5</position>
<output>
<ID>OUT_0</ID>7 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>417</ID>
<type>AA_LABEL</type>
<position>124,-223</position>
<gparam>LABEL_TEXT borrow=a'b</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>28</ID>
<type>AA_TOGGLE</type>
<position>52,-15.5</position>
<output>
<ID>OUT_0</ID>8 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>418</ID>
<type>AA_LABEL</type>
<position>6.5,-289.5</position>
<gparam>LABEL_TEXT Full Adder</gparam>
<gparam>TEXT_HEIGHT 7</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>29</ID>
<type>AA_TOGGLE</type>
<position>23,-7.5</position>
<output>
<ID>OUT_0</ID>9 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>30</ID>
<type>AA_TOGGLE</type>
<position>23,-9.5</position>
<output>
<ID>OUT_0</ID>10 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>420</ID>
<type>AI_XOR3</type>
<position>41,-263.5</position>
<input>
<ID>IN_0</ID>229 </input>
<input>
<ID>IN_1</ID>230 </input>
<input>
<ID>IN_2</ID>231 </input>
<output>
<ID>OUT</ID>232 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>31</ID>
<type>AA_TOGGLE</type>
<position>23,-3</position>
<output>
<ID>OUT_0</ID>11 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>422</ID>
<type>AA_AND2</type>
<position>47,-274.5</position>
<input>
<ID>IN_0</ID>229 </input>
<input>
<ID>IN_1</ID>230 </input>
<output>
<ID>OUT</ID>226 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>33</ID>
<type>GA_LED</type>
<position>34.5,-3</position>
<input>
<ID>N_in0</ID>12 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>423</ID>
<type>AA_AND2</type>
<position>47,-280.5</position>
<input>
<ID>IN_0</ID>230 </input>
<input>
<ID>IN_1</ID>231 </input>
<output>
<ID>OUT</ID>227 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>34</ID>
<type>GA_LED</type>
<position>65,-9</position>
<input>
<ID>N_in0</ID>14 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>424</ID>
<type>AA_AND2</type>
<position>47,-286</position>
<input>
<ID>IN_0</ID>229 </input>
<input>
<ID>IN_1</ID>231 </input>
<output>
<ID>OUT</ID>228 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>35</ID>
<type>GA_LED</type>
<position>34.5,-8.5</position>
<input>
<ID>N_in0</ID>13 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>36</ID>
<type>GA_LED</type>
<position>65,-14.5</position>
<input>
<ID>N_in0</ID>16 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>426</ID>
<type>AE_OR3</type>
<position>59,-280.5</position>
<input>
<ID>IN_0</ID>226 </input>
<input>
<ID>IN_1</ID>227 </input>
<input>
<ID>IN_2</ID>228 </input>
<output>
<ID>OUT</ID>233 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>37</ID>
<type>AA_LABEL</type>
<position>21,-2.5</position>
<gparam>LABEL_TEXT a</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>38</ID>
<type>AA_LABEL</type>
<position>21,-7</position>
<gparam>LABEL_TEXT a</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>428</ID>
<type>AA_TOGGLE</type>
<position>24.5,-258</position>
<output>
<ID>OUT_0</ID>229 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>39</ID>
<type>AA_LABEL</type>
<position>50,-13</position>
<gparam>LABEL_TEXT a</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>429</ID>
<type>AA_TOGGLE</type>
<position>28,-258</position>
<output>
<ID>OUT_0</ID>230 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>40</ID>
<type>AA_LABEL</type>
<position>50,-7.5</position>
<gparam>LABEL_TEXT a</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>430</ID>
<type>AA_TOGGLE</type>
<position>31.5,-258</position>
<output>
<ID>OUT_0</ID>231 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>41</ID>
<type>AA_LABEL</type>
<position>21,-9.5</position>
<gparam>LABEL_TEXT b</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>42</ID>
<type>AA_LABEL</type>
<position>50,-15.5</position>
<gparam>LABEL_TEXT b</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>432</ID>
<type>GA_LED</type>
<position>48,-264</position>
<input>
<ID>N_in0</ID>232 </input>
<input>
<ID>N_in3</ID>232 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>43</ID>
<type>AA_LABEL</type>
<position>50,-9.5</position>
<gparam>LABEL_TEXT b</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>433</ID>
<type>GA_LED</type>
<position>65.5,-280.5</position>
<input>
<ID>N_in0</ID>233 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>44</ID>
<type>AA_LABEL</type>
<position>70,-14</position>
<gparam>LABEL_TEXT y=(a.b)'</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>45</ID>
<type>AA_LABEL</type>
<position>38.5,-8</position>
<gparam>LABEL_TEXT y=a+b</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>435</ID>
<type>AA_LABEL</type>
<position>31.5,-255.5</position>
<gparam>LABEL_TEXT cin</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>46</ID>
<type>AA_LABEL</type>
<position>70,-8.5</position>
<gparam>LABEL_TEXT y=(a+b)'</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>47</ID>
<type>AA_LABEL</type>
<position>38,-2.5</position>
<gparam>LABEL_TEXT y=a'</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>437</ID>
<type>AA_LABEL</type>
<position>48,-261</position>
<gparam>LABEL_TEXT sum</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>438</ID>
<type>AA_LABEL</type>
<position>65.5,-278</position>
<gparam>LABEL_TEXT carry</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>439</ID>
<type>AA_LABEL</type>
<position>24,-255.5</position>
<gparam>LABEL_TEXT a</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>440</ID>
<type>AA_LABEL</type>
<position>28,-255.5</position>
<gparam>LABEL_TEXT b</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>51</ID>
<type>AA_LABEL</type>
<position>10,-35</position>
<gparam>LABEL_TEXT NAND as universal</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>53</ID>
<type>BA_NAND2</type>
<position>23.5,-23.5</position>
<input>
<ID>IN_0</ID>17 </input>
<input>
<ID>IN_1</ID>17 </input>
<output>
<ID>OUT</ID>18 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>55</ID>
<type>AA_TOGGLE</type>
<position>17,-23.5</position>
<output>
<ID>OUT_0</ID>17 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>445</ID>
<type>AA_AND3</type>
<position>140,-267</position>
<input>
<ID>IN_0</ID>246 </input>
<input>
<ID>IN_1</ID>247 </input>
<input>
<ID>IN_2</ID>248 </input>
<output>
<ID>OUT</ID>235 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>446</ID>
<type>AA_AND3</type>
<position>141,-275.5</position>
<input>
<ID>IN_0</ID>246 </input>
<input>
<ID>IN_1</ID>244 </input>
<input>
<ID>IN_2</ID>249 </input>
<output>
<ID>OUT</ID>236 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>57</ID>
<type>GA_LED</type>
<position>28.5,-23.5</position>
<input>
<ID>N_in0</ID>18 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>447</ID>
<type>AA_AND3</type>
<position>140,-284.5</position>
<input>
<ID>IN_0</ID>250 </input>
<input>
<ID>IN_1</ID>247 </input>
<input>
<ID>IN_2</ID>249 </input>
<output>
<ID>OUT</ID>237 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>448</ID>
<type>AA_AND3</type>
<position>140,-294</position>
<input>
<ID>IN_0</ID>250 </input>
<input>
<ID>IN_1</ID>244 </input>
<input>
<ID>IN_2</ID>248 </input>
<output>
<ID>OUT</ID>238 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>59</ID>
<type>BA_NAND2</type>
<position>41,-24</position>
<input>
<ID>IN_0</ID>20 </input>
<input>
<ID>IN_1</ID>21 </input>
<output>
<ID>OUT</ID>19 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>449</ID>
<type>AA_AND3</type>
<position>140,-308.5</position>
<input>
<ID>IN_0</ID>250 </input>
<input>
<ID>IN_1</ID>247 </input>
<input>
<ID>IN_2</ID>248 </input>
<output>
<ID>OUT</ID>239 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>450</ID>
<type>AA_AND3</type>
<position>140,-318</position>
<input>
<ID>IN_0</ID>246 </input>
<input>
<ID>IN_1</ID>244 </input>
<input>
<ID>IN_2</ID>248 </input>
<output>
<ID>OUT</ID>240 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>61</ID>
<type>BA_NAND2</type>
<position>49.5,-24</position>
<input>
<ID>IN_0</ID>19 </input>
<input>
<ID>IN_1</ID>19 </input>
<output>
<ID>OUT</ID>22 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>451</ID>
<type>AA_AND3</type>
<position>140,-327</position>
<input>
<ID>IN_0</ID>250 </input>
<input>
<ID>IN_1</ID>244 </input>
<input>
<ID>IN_2</ID>249 </input>
<output>
<ID>OUT</ID>241 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>62</ID>
<type>AA_TOGGLE</type>
<position>36,-23</position>
<output>
<ID>OUT_0</ID>20 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>452</ID>
<type>AA_AND3</type>
<position>140,-336.5</position>
<output>
<ID>OUT</ID>242 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>63</ID>
<type>AA_TOGGLE</type>
<position>36,-25</position>
<output>
<ID>OUT_0</ID>21 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>64</ID>
<type>GA_LED</type>
<position>54.5,-24</position>
<input>
<ID>N_in0</ID>22 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>454</ID>
<type>AE_SMALL_INVERTER</type>
<position>33.5,-171.5</position>
<input>
<ID>IN_0</ID>195 </input>
<output>
<ID>OUT_0</ID>234 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>66</ID>
<type>BA_NAND2</type>
<position>72.5,-23.5</position>
<input>
<ID>IN_0</ID>26 </input>
<input>
<ID>IN_1</ID>26 </input>
<output>
<ID>OUT</ID>23 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>456</ID>
<type>AA_TOGGLE</type>
<position>99,-251</position>
<output>
<ID>OUT_0</ID>250 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>457</ID>
<type>AA_TOGGLE</type>
<position>111,-251</position>
<output>
<ID>OUT_0</ID>244 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>68</ID>
<type>BA_NAND2</type>
<position>72.5,-29</position>
<input>
<ID>IN_0</ID>27 </input>
<input>
<ID>IN_1</ID>27 </input>
<output>
<ID>OUT</ID>24 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>458</ID>
<type>AA_TOGGLE</type>
<position>122.5,-251</position>
<output>
<ID>OUT_0</ID>248 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>70</ID>
<type>BA_NAND2</type>
<position>81,-26.5</position>
<input>
<ID>IN_0</ID>23 </input>
<input>
<ID>IN_1</ID>24 </input>
<output>
<ID>OUT</ID>28 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>460</ID>
<type>AE_SMALL_INVERTER</type>
<position>103,-257</position>
<input>
<ID>IN_0</ID>250 </input>
<output>
<ID>OUT_0</ID>246 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>71</ID>
<type>AA_TOGGLE</type>
<position>65,-23.5</position>
<output>
<ID>OUT_0</ID>26 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>461</ID>
<type>AE_SMALL_INVERTER</type>
<position>116,-257</position>
<input>
<ID>IN_0</ID>244 </input>
<output>
<ID>OUT_0</ID>247 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>72</ID>
<type>AA_TOGGLE</type>
<position>65,-29</position>
<output>
<ID>OUT_0</ID>27 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>462</ID>
<type>AE_SMALL_INVERTER</type>
<position>128,-257</position>
<input>
<ID>IN_0</ID>248 </input>
<output>
<ID>OUT_0</ID>249 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>73</ID>
<type>AA_TOGGLE</type>
<position>18,-35.5</position>
<output>
<ID>OUT_0</ID>36 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>74</ID>
<type>GA_LED</type>
<position>86,-26.5</position>
<input>
<ID>N_in0</ID>28 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>464</ID>
<type>AE_OR4</type>
<position>165,-282</position>
<input>
<ID>IN_0</ID>235 </input>
<input>
<ID>IN_1</ID>236 </input>
<input>
<ID>IN_2</ID>237 </input>
<input>
<ID>IN_3</ID>238 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>465</ID>
<type>AE_OR4</type>
<position>164,-321.5</position>
<input>
<ID>IN_0</ID>239 </input>
<input>
<ID>IN_1</ID>240 </input>
<input>
<ID>IN_2</ID>241 </input>
<input>
<ID>IN_3</ID>242 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>76</ID>
<type>BA_NAND2</type>
<position>25.5,-39.5</position>
<input>
<ID>IN_0</ID>36 </input>
<input>
<ID>IN_1</ID>35 </input>
<output>
<ID>OUT</ID>34 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>77</ID>
<type>BA_NAND2</type>
<position>33.5,-36.5</position>
<input>
<ID>IN_0</ID>36 </input>
<input>
<ID>IN_1</ID>34 </input>
<output>
<ID>OUT</ID>31 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>78</ID>
<type>BA_NAND2</type>
<position>33,-43</position>
<input>
<ID>IN_0</ID>34 </input>
<input>
<ID>IN_1</ID>35 </input>
<output>
<ID>OUT</ID>32 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>79</ID>
<type>BA_NAND2</type>
<position>42,-40</position>
<input>
<ID>IN_0</ID>31 </input>
<input>
<ID>IN_1</ID>32 </input>
<output>
<ID>OUT</ID>37 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>80</ID>
<type>BA_NAND2</type>
<position>82,-37</position>
<input>
<ID>IN_0</ID>42 </input>
<input>
<ID>IN_1</ID>45 </input>
<output>
<ID>OUT</ID>38 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>81</ID>
<type>BA_NAND2</type>
<position>82.5,-43</position>
<input>
<ID>IN_0</ID>42 </input>
<input>
<ID>IN_1</ID>42 </input>
<output>
<ID>OUT</ID>40 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>82</ID>
<type>BA_NAND2</type>
<position>91.5,-45.5</position>
<input>
<ID>IN_0</ID>40 </input>
<input>
<ID>IN_1</ID>41 </input>
<output>
<ID>OUT</ID>39 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>83</ID>
<type>BA_NAND2</type>
<position>101.5,-42.5</position>
<input>
<ID>IN_0</ID>38 </input>
<input>
<ID>IN_1</ID>39 </input>
<output>
<ID>OUT</ID>46 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>84</ID>
<type>BA_NAND2</type>
<position>82,-48</position>
<input>
<ID>IN_0</ID>45 </input>
<input>
<ID>IN_1</ID>45 </input>
<output>
<ID>OUT</ID>41 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>85</ID>
<type>AA_TOGGLE</type>
<position>18,-42.5</position>
<output>
<ID>OUT_0</ID>35 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>87</ID>
<type>GA_LED</type>
<position>48,-40</position>
<input>
<ID>N_in0</ID>37 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>89</ID>
<type>AA_TOGGLE</type>
<position>71.5,-36</position>
<output>
<ID>OUT_0</ID>42 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>90</ID>
<type>AA_TOGGLE</type>
<position>71.5,-38</position>
<output>
<ID>OUT_0</ID>45 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>91</ID>
<type>AA_LABEL</type>
<position>69.5,-35.5</position>
<gparam>LABEL_TEXT a</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>92</ID>
<type>AA_LABEL</type>
<position>69.5,-37.5</position>
<gparam>LABEL_TEXT b</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>97</ID>
<type>GA_LED</type>
<position>106.5,-42.5</position>
<input>
<ID>N_in0</ID>46 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>101</ID>
<type>AA_TOGGLE</type>
<position>84.5,-10.5</position>
<output>
<ID>OUT_0</ID>51 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>102</ID>
<type>AA_TOGGLE</type>
<position>84.5,-8.5</position>
<output>
<ID>OUT_0</ID>50 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>103</ID>
<type>GA_LED</type>
<position>97.5,-9.5</position>
<input>
<ID>N_in0</ID>52 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>104</ID>
<type>AA_LABEL</type>
<position>82.5,-8</position>
<gparam>LABEL_TEXT a</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>105</ID>
<type>AA_LABEL</type>
<position>82.5,-10</position>
<gparam>LABEL_TEXT b</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>106</ID>
<type>AA_LABEL</type>
<position>103,-9</position>
<gparam>LABEL_TEXT y=ab'+a'b</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>110</ID>
<type>AI_XOR2</type>
<position>92,-9.5</position>
<input>
<ID>IN_0</ID>50 </input>
<input>
<ID>IN_1</ID>51 </input>
<output>
<ID>OUT</ID>52 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>112</ID>
<type>AO_XNOR2</type>
<position>92.5,-15</position>
<input>
<ID>IN_0</ID>56 </input>
<input>
<ID>IN_1</ID>63 </input>
<output>
<ID>OUT</ID>65 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>113</ID>
<type>AA_TOGGLE</type>
<position>84.5,-16</position>
<output>
<ID>OUT_0</ID>63 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>114</ID>
<type>AA_TOGGLE</type>
<position>84.5,-13.5</position>
<output>
<ID>OUT_0</ID>56 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>115</ID>
<type>GA_LED</type>
<position>98,-15</position>
<input>
<ID>N_in0</ID>65 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>116</ID>
<type>AA_LABEL</type>
<position>82.5,-13</position>
<gparam>LABEL_TEXT a</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>117</ID>
<type>AA_LABEL</type>
<position>82.5,-15.5</position>
<gparam>LABEL_TEXT b</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>118</ID>
<type>AA_LABEL</type>
<position>103.5,-14.5</position>
<gparam>LABEL_TEXT y=ab+a'b'</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>127</ID>
<type>AA_LABEL</type>
<position>9,-68.5</position>
<gparam>LABEL_TEXT NOR as universal</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>128</ID>
<type>AA_LABEL</type>
<position>15,-23</position>
<gparam>LABEL_TEXT a</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>129</ID>
<type>AA_LABEL</type>
<position>16,-35</position>
<gparam>LABEL_TEXT a</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>130</ID>
<type>AA_LABEL</type>
<position>34,-22.5</position>
<gparam>LABEL_TEXT a</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>131</ID>
<type>AA_LABEL</type>
<position>63,-23</position>
<gparam>LABEL_TEXT a</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>132</ID>
<type>AA_LABEL</type>
<position>16,-42</position>
<gparam>LABEL_TEXT b</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>133</ID>
<type>AA_LABEL</type>
<position>34,-25</position>
<gparam>LABEL_TEXT b</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>134</ID>
<type>AA_LABEL</type>
<position>63,-29</position>
<gparam>LABEL_TEXT b</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>136</ID>
<type>AA_TOGGLE</type>
<position>19.5,-59</position>
<output>
<ID>OUT_0</ID>90 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>137</ID>
<type>GA_LED</type>
<position>31,-59</position>
<input>
<ID>N_in0</ID>91 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>140</ID>
<type>AA_TOGGLE</type>
<position>38.5,-58.5</position>
<output>
<ID>OUT_0</ID>94 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>141</ID>
<type>AA_TOGGLE</type>
<position>38.5,-60.5</position>
<output>
<ID>OUT_0</ID>95 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>142</ID>
<type>GA_LED</type>
<position>57,-59.5</position>
<input>
<ID>N_in0</ID>93 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>146</ID>
<type>AA_TOGGLE</type>
<position>67.5,-59</position>
<output>
<ID>OUT_0</ID>96 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>147</ID>
<type>AA_TOGGLE</type>
<position>67.5,-64.5</position>
<output>
<ID>OUT_0</ID>97 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>148</ID>
<type>AA_TOGGLE</type>
<position>20.5,-71</position>
<output>
<ID>OUT_0</ID>81 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>149</ID>
<type>GA_LED</type>
<position>88.5,-62</position>
<input>
<ID>N_in0</ID>100 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>159</ID>
<type>AA_TOGGLE</type>
<position>20.5,-79</position>
<output>
<ID>OUT_0</ID>80 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>160</ID>
<type>GA_LED</type>
<position>50.5,-75.5</position>
<input>
<ID>N_in0</ID>103 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>166</ID>
<type>AA_LABEL</type>
<position>17.5,-58.5</position>
<gparam>LABEL_TEXT a</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>167</ID>
<type>AA_LABEL</type>
<position>18.5,-70.5</position>
<gparam>LABEL_TEXT a</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>168</ID>
<type>AA_LABEL</type>
<position>36.5,-58</position>
<gparam>LABEL_TEXT a</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>169</ID>
<type>AA_LABEL</type>
<position>65.5,-58.5</position>
<gparam>LABEL_TEXT a</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>170</ID>
<type>AA_LABEL</type>
<position>18.5,-77.5</position>
<gparam>LABEL_TEXT b</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>171</ID>
<type>AA_LABEL</type>
<position>36.5,-60.5</position>
<gparam>LABEL_TEXT b</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>172</ID>
<type>AA_LABEL</type>
<position>65.5,-64.5</position>
<gparam>LABEL_TEXT b</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>174</ID>
<type>BE_NOR2</type>
<position>26,-59</position>
<input>
<ID>IN_0</ID>90 </input>
<input>
<ID>IN_1</ID>90 </input>
<output>
<ID>OUT</ID>91 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>175</ID>
<type>BE_NOR2</type>
<position>45,-59.5</position>
<input>
<ID>IN_0</ID>94 </input>
<input>
<ID>IN_1</ID>95 </input>
<output>
<ID>OUT</ID>92 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>176</ID>
<type>BE_NOR2</type>
<position>52,-59.5</position>
<input>
<ID>IN_0</ID>92 </input>
<input>
<ID>IN_1</ID>92 </input>
<output>
<ID>OUT</ID>93 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>177</ID>
<type>BE_NOR2</type>
<position>75,-58.5</position>
<input>
<ID>IN_0</ID>96 </input>
<input>
<ID>IN_1</ID>96 </input>
<output>
<ID>OUT</ID>98 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>178</ID>
<type>BE_NOR2</type>
<position>75,-64.5</position>
<input>
<ID>IN_0</ID>97 </input>
<input>
<ID>IN_1</ID>97 </input>
<output>
<ID>OUT</ID>99 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>179</ID>
<type>BE_NOR2</type>
<position>83.5,-62</position>
<input>
<ID>IN_0</ID>98 </input>
<input>
<ID>IN_1</ID>99 </input>
<output>
<ID>OUT</ID>100 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>180</ID>
<type>BE_NOR2</type>
<position>28.5,-75</position>
<input>
<ID>IN_0</ID>81 </input>
<input>
<ID>IN_1</ID>80 </input>
<output>
<ID>OUT</ID>79 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>181</ID>
<type>BE_NOR2</type>
<position>38,-72</position>
<input>
<ID>IN_0</ID>81 </input>
<input>
<ID>IN_1</ID>79 </input>
<output>
<ID>OUT</ID>101 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>182</ID>
<type>BE_NOR2</type>
<position>37.5,-78</position>
<input>
<ID>IN_0</ID>79 </input>
<input>
<ID>IN_1</ID>80 </input>
<output>
<ID>OUT</ID>102 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>183</ID>
<type>BE_NOR2</type>
<position>45.5,-75.5</position>
<input>
<ID>IN_0</ID>101 </input>
<input>
<ID>IN_1</ID>102 </input>
<output>
<ID>OUT</ID>103 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>193</ID>
<type>AA_TOGGLE</type>
<position>63.5,-72.5</position>
<output>
<ID>OUT_0</ID>112 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>194</ID>
<type>AA_TOGGLE</type>
<position>63.5,-80.5</position>
<output>
<ID>OUT_0</ID>111 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>195</ID>
<type>GA_LED</type>
<position>102,-77</position>
<input>
<ID>N_in0</ID>117 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>196</ID>
<type>AA_LABEL</type>
<position>61.5,-72</position>
<gparam>LABEL_TEXT a</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>197</ID>
<type>AA_LABEL</type>
<position>61.5,-79</position>
<gparam>LABEL_TEXT b</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>198</ID>
<type>BE_NOR2</type>
<position>71.5,-76.5</position>
<input>
<ID>IN_0</ID>112 </input>
<input>
<ID>IN_1</ID>111 </input>
<output>
<ID>OUT</ID>110 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>199</ID>
<type>BE_NOR2</type>
<position>81,-73.5</position>
<input>
<ID>IN_0</ID>112 </input>
<input>
<ID>IN_1</ID>110 </input>
<output>
<ID>OUT</ID>113 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>200</ID>
<type>BE_NOR2</type>
<position>80.5,-79.5</position>
<input>
<ID>IN_0</ID>110 </input>
<input>
<ID>IN_1</ID>111 </input>
<output>
<ID>OUT</ID>114 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>201</ID>
<type>BE_NOR2</type>
<position>88.5,-77</position>
<input>
<ID>IN_0</ID>113 </input>
<input>
<ID>IN_1</ID>114 </input>
<output>
<ID>OUT</ID>116 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>202</ID>
<type>BE_NOR2</type>
<position>96.5,-77</position>
<input>
<ID>IN_0</ID>116 </input>
<input>
<ID>IN_1</ID>116 </input>
<output>
<ID>OUT</ID>117 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>203</ID>
<type>AA_LABEL</type>
<position>28.5,-20.5</position>
<gparam>LABEL_TEXT y=a'</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>204</ID>
<type>AA_LABEL</type>
<position>31,-56.5</position>
<gparam>LABEL_TEXT y=a'</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>205</ID>
<type>AA_LABEL</type>
<position>55,-21</position>
<gparam>LABEL_TEXT y=a.b</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>206</ID>
<type>AA_LABEL</type>
<position>89,-59</position>
<gparam>LABEL_TEXT y=a.b</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>207</ID>
<type>AA_LABEL</type>
<position>87,-23.5</position>
<gparam>LABEL_TEXT y=a+b</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>208</ID>
<type>AA_LABEL</type>
<position>57,-57</position>
<gparam>LABEL_TEXT y=a+b</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>209</ID>
<type>AA_LABEL</type>
<position>54,-39.5</position>
<gparam>LABEL_TEXT y=ab'+a'b</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>210</ID>
<type>AA_LABEL</type>
<position>108,-76.5</position>
<gparam>LABEL_TEXT y=ab'+a'b</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>211</ID>
<type>AA_LABEL</type>
<position>112.5,-42</position>
<gparam>LABEL_TEXT y=ab+a'b'</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>212</ID>
<type>AA_LABEL</type>
<position>52,-73</position>
<gparam>LABEL_TEXT y=ab+a'b'</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>213</ID>
<type>AA_LABEL</type>
<position>9,-119.5</position>
<gparam>LABEL_TEXT Half Adder</gparam>
<gparam>TEXT_HEIGHT 7</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>215</ID>
<type>AI_XOR2</type>
<position>31,-96.5</position>
<input>
<ID>IN_0</ID>118 </input>
<input>
<ID>IN_1</ID>119 </input>
<output>
<ID>OUT</ID>120 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>217</ID>
<type>AA_AND2</type>
<position>31,-103.5</position>
<input>
<ID>IN_0</ID>118 </input>
<input>
<ID>IN_1</ID>119 </input>
<output>
<ID>OUT</ID>122 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>218</ID>
<type>AA_TOGGLE</type>
<position>21.5,-95.5</position>
<output>
<ID>OUT_0</ID>118 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>219</ID>
<type>AA_LABEL</type>
<position>19.5,-95</position>
<gparam>LABEL_TEXT a</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>220</ID>
<type>AA_TOGGLE</type>
<position>21.5,-98.5</position>
<output>
<ID>OUT_0</ID>119 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>221</ID>
<type>AA_LABEL</type>
<position>19.5,-98</position>
<gparam>LABEL_TEXT b</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>223</ID>
<type>GA_LED</type>
<position>37.5,-96.5</position>
<input>
<ID>N_in0</ID>120 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>225</ID>
<type>GA_LED</type>
<position>37.5,-103.5</position>
<input>
<ID>N_in0</ID>122 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>227</ID>
<type>AA_TOGGLE</type>
<position>63.5,-91.5</position>
<output>
<ID>OUT_0</ID>123 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>228</ID>
<type>AA_TOGGLE</type>
<position>74,-91</position>
<output>
<ID>OUT_0</ID>124 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>230</ID>
<type>AE_SMALL_INVERTER</type>
<position>68.5,-96.5</position>
<input>
<ID>IN_0</ID>123 </input>
<output>
<ID>OUT_0</ID>127 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>232</ID>
<type>AE_SMALL_INVERTER</type>
<position>79,-96</position>
<input>
<ID>IN_0</ID>124 </input>
<output>
<ID>OUT_0</ID>128 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>234</ID>
<type>AA_AND2</type>
<position>89,-101</position>
<input>
<ID>IN_0</ID>123 </input>
<input>
<ID>IN_1</ID>128 </input>
<output>
<ID>OUT</ID>125 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>235</ID>
<type>AA_AND2</type>
<position>89,-107</position>
<input>
<ID>IN_0</ID>127 </input>
<input>
<ID>IN_1</ID>124 </input>
<output>
<ID>OUT</ID>126 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>236</ID>
<type>AA_AND2</type>
<position>93,-112</position>
<input>
<ID>IN_0</ID>123 </input>
<input>
<ID>IN_1</ID>124 </input>
<output>
<ID>OUT</ID>130 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>238</ID>
<type>AE_OR2</type>
<position>98.5,-104</position>
<input>
<ID>IN_0</ID>125 </input>
<input>
<ID>IN_1</ID>126 </input>
<output>
<ID>OUT</ID>129 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>240</ID>
<type>GA_LED</type>
<position>106.5,-104</position>
<input>
<ID>N_in0</ID>129 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>242</ID>
<type>GA_LED</type>
<position>101,-114</position>
<input>
<ID>N_in0</ID>130 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>244</ID>
<type>AA_LABEL</type>
<position>39,-94</position>
<gparam>LABEL_TEXT sum=ab'+a'b</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>245</ID>
<type>AA_LABEL</type>
<position>107,-101</position>
<gparam>LABEL_TEXT sum=ab'+a'b</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>247</ID>
<type>AA_LABEL</type>
<position>37.5,-100.5</position>
<gparam>LABEL_TEXT carry=ab</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>248</ID>
<type>AA_LABEL</type>
<position>101,-111.5</position>
<gparam>LABEL_TEXT carry=ab</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>250</ID>
<type>AA_LABEL</type>
<position>10,-7.5</position>
<gparam>LABEL_TEXT Basic Gates</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>251</ID>
<type>AA_LABEL</type>
<position>63.5,-89</position>
<gparam>LABEL_TEXT a</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>254</ID>
<type>AA_LABEL</type>
<position>74,-88.5</position>
<gparam>LABEL_TEXT b</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>296</ID>
<type>AA_TOGGLE</type>
<position>17.5,-122</position>
<output>
<ID>OUT_0</ID>156 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>297</ID>
<type>AA_LABEL</type>
<position>17.5,-119.5</position>
<gparam>LABEL_TEXT a</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>298</ID>
<type>AA_LABEL</type>
<position>27.5,-119.5</position>
<gparam>LABEL_TEXT b</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>299</ID>
<type>BA_NAND2</type>
<position>23,-127.5</position>
<input>
<ID>IN_0</ID>156 </input>
<input>
<ID>IN_1</ID>156 </input>
<output>
<ID>OUT</ID>157 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>300</ID>
<type>AA_TOGGLE</type>
<position>27.5,-122</position>
<output>
<ID>OUT_0</ID>152 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>301</ID>
<type>BA_NAND2</type>
<position>32.5,-127</position>
<input>
<ID>IN_0</ID>152 </input>
<input>
<ID>IN_1</ID>152 </input>
<output>
<ID>OUT</ID>158 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>302</ID>
<type>BA_NAND2</type>
<position>45,-134</position>
<input>
<ID>IN_0</ID>156 </input>
<input>
<ID>IN_1</ID>158 </input>
<output>
<ID>OUT</ID>153 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>303</ID>
<type>BA_NAND2</type>
<position>45,-139</position>
<input>
<ID>IN_0</ID>157 </input>
<input>
<ID>IN_1</ID>152 </input>
<output>
<ID>OUT</ID>154 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>304</ID>
<type>BA_NAND2</type>
<position>45.5,-147</position>
<input>
<ID>IN_0</ID>156 </input>
<input>
<ID>IN_1</ID>152 </input>
<output>
<ID>OUT</ID>155 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>305</ID>
<type>BA_NAND2</type>
<position>56.5,-147</position>
<input>
<ID>IN_0</ID>155 </input>
<input>
<ID>IN_1</ID>155 </input>
<output>
<ID>OUT</ID>160 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>306</ID>
<type>BA_NAND2</type>
<position>56.5,-136.5</position>
<input>
<ID>IN_0</ID>153 </input>
<input>
<ID>IN_1</ID>154 </input>
<output>
<ID>OUT</ID>159 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>307</ID>
<type>GA_LED</type>
<position>63.5,-136.5</position>
<input>
<ID>N_in0</ID>159 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>308</ID>
<type>GA_LED</type>
<position>64,-147</position>
<input>
<ID>N_in0</ID>160 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>309</ID>
<type>AA_LABEL</type>
<position>64.5,-134</position>
<gparam>LABEL_TEXT sum=ab'+a'b</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>310</ID>
<type>AA_LABEL</type>
<position>64,-144</position>
<gparam>LABEL_TEXT carry=ab</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>311</ID>
<type>AA_TOGGLE</type>
<position>77,-124.5</position>
<output>
<ID>OUT_0</ID>185 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>312</ID>
<type>AA_LABEL</type>
<position>77,-122</position>
<gparam>LABEL_TEXT a</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>313</ID>
<type>AA_LABEL</type>
<position>87,-122</position>
<gparam>LABEL_TEXT b</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>327</ID>
<type>BE_NOR2</type>
<position>104.5,-136</position>
<input>
<ID>IN_0</ID>181 </input>
<input>
<ID>IN_1</ID>183 </input>
<output>
<ID>OUT</ID>186 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>343</ID>
<type>BE_NOR2</type>
<position>104.5,-141</position>
<input>
<ID>IN_0</ID>185 </input>
<input>
<ID>IN_1</ID>184 </input>
<output>
<ID>OUT</ID>187 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>344</ID>
<type>BE_NOR2</type>
<position>104,-150</position>
<input>
<ID>IN_0</ID>181 </input>
<input>
<ID>IN_1</ID>184 </input>
<output>
<ID>OUT</ID>188 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>345</ID>
<type>BE_NOR2</type>
<position>114.5,-138.5</position>
<input>
<ID>IN_0</ID>186 </input>
<input>
<ID>IN_1</ID>187 </input>
<output>
<ID>OUT</ID>190 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>347</ID>
<type>BE_NOR2</type>
<position>81.5,-131.5</position>
<input>
<ID>IN_0</ID>185 </input>
<input>
<ID>IN_1</ID>185 </input>
<output>
<ID>OUT</ID>181 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>348</ID>
<type>AA_TOGGLE</type>
<position>87,-124.5</position>
<output>
<ID>OUT_0</ID>183 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>349</ID>
<type>BE_NOR2</type>
<position>91,-131.5</position>
<input>
<ID>IN_0</ID>183 </input>
<input>
<ID>IN_1</ID>183 </input>
<output>
<ID>OUT</ID>184 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>350</ID>
<type>GA_LED</type>
<position>129.5,-138.5</position>
<input>
<ID>N_in0</ID>189 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>351</ID>
<type>GA_LED</type>
<position>112,-150</position>
<input>
<ID>N_in0</ID>188 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>352</ID>
<type>AA_LABEL</type>
<position>111.5,-147.5</position>
<gparam>LABEL_TEXT carry=ab</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>353</ID>
<type>BE_NOR2</type>
<position>123,-138.5</position>
<input>
<ID>IN_0</ID>190 </input>
<input>
<ID>IN_1</ID>190 </input>
<output>
<ID>OUT</ID>189 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>354</ID>
<type>AA_LABEL</type>
<position>131,-135.5</position>
<gparam>LABEL_TEXT sum=ab'+a'b</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>355</ID>
<type>AA_LABEL</type>
<position>7.5,-200.5</position>
<gparam>LABEL_TEXT Half subtractor</gparam>
<gparam>TEXT_HEIGHT 7</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>356</ID>
<type>AI_XOR2</type>
<position>37,-167.5</position>
<input>
<ID>IN_0</ID>195 </input>
<input>
<ID>IN_1</ID>192 </input>
<output>
<ID>OUT</ID>193 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>357</ID>
<type>AA_AND2</type>
<position>37,-174.5</position>
<input>
<ID>IN_0</ID>234 </input>
<input>
<ID>IN_1</ID>192 </input>
<output>
<ID>OUT</ID>194 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>358</ID>
<type>AA_TOGGLE</type>
<position>27.5,-166.5</position>
<output>
<ID>OUT_0</ID>195 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>359</ID>
<type>AA_LABEL</type>
<position>25.5,-166</position>
<gparam>LABEL_TEXT a</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>360</ID>
<type>AA_TOGGLE</type>
<position>27.5,-169.5</position>
<output>
<ID>OUT_0</ID>192 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>361</ID>
<type>AA_LABEL</type>
<position>25.5,-169</position>
<gparam>LABEL_TEXT b</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>362</ID>
<type>GA_LED</type>
<position>43.5,-167.5</position>
<input>
<ID>N_in0</ID>193 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>363</ID>
<type>GA_LED</type>
<position>43.5,-174.5</position>
<input>
<ID>N_in0</ID>194 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>364</ID>
<type>AA_LABEL</type>
<position>44.5,-165</position>
<gparam>LABEL_TEXT diff=ab'+a'b</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>365</ID>
<type>AA_LABEL</type>
<position>43.5,-171.5</position>
<gparam>LABEL_TEXT borrow=a'b</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>368</ID>
<type>AA_TOGGLE</type>
<position>78,-164</position>
<output>
<ID>OUT_0</ID>205 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>369</ID>
<type>AA_TOGGLE</type>
<position>88.5,-163.5</position>
<output>
<ID>OUT_0</ID>198 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>370</ID>
<type>AE_SMALL_INVERTER</type>
<position>83,-169</position>
<input>
<ID>IN_0</ID>205 </input>
<output>
<ID>OUT_0</ID>201 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>371</ID>
<type>AE_SMALL_INVERTER</type>
<position>93.5,-168.5</position>
<input>
<ID>IN_0</ID>198 </input>
<output>
<ID>OUT_0</ID>202 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>372</ID>
<type>AA_AND2</type>
<position>103.5,-173.5</position>
<input>
<ID>IN_0</ID>205 </input>
<input>
<ID>IN_1</ID>202 </input>
<output>
<ID>OUT</ID>199 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>373</ID>
<type>AA_AND2</type>
<position>103.5,-179.5</position>
<input>
<ID>IN_0</ID>201 </input>
<input>
<ID>IN_1</ID>198 </input>
<output>
<ID>OUT</ID>200 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>374</ID>
<type>AA_AND2</type>
<position>107.5,-184.5</position>
<input>
<ID>IN_0</ID>201 </input>
<input>
<ID>IN_1</ID>198 </input>
<output>
<ID>OUT</ID>204 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>375</ID>
<type>AE_OR2</type>
<position>113,-176.5</position>
<input>
<ID>IN_0</ID>199 </input>
<input>
<ID>IN_1</ID>200 </input>
<output>
<ID>OUT</ID>203 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>376</ID>
<type>GA_LED</type>
<position>121,-176.5</position>
<input>
<ID>N_in0</ID>203 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>377</ID>
<type>GA_LED</type>
<position>115.5,-186.5</position>
<input>
<ID>N_in0</ID>204 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>380</ID>
<type>AA_LABEL</type>
<position>78,-161.5</position>
<gparam>LABEL_TEXT a</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>381</ID>
<type>AA_LABEL</type>
<position>88.5,-161</position>
<gparam>LABEL_TEXT b</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>382</ID>
<type>AA_LABEL</type>
<position>121.5,-173.5</position>
<gparam>LABEL_TEXT diff=ab'+a'b</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>383</ID>
<type>AA_LABEL</type>
<position>117.5,-182.5</position>
<gparam>LABEL_TEXT borrow=a'b</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>384</ID>
<type>AA_TOGGLE</type>
<position>23.5,-200</position>
<output>
<ID>OUT_0</ID>215 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>385</ID>
<type>AA_LABEL</type>
<position>23.5,-197.5</position>
<gparam>LABEL_TEXT a</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>386</ID>
<type>AA_LABEL</type>
<position>33.5,-197.5</position>
<gparam>LABEL_TEXT b</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>387</ID>
<type>BA_NAND2</type>
<position>29,-206</position>
<input>
<ID>IN_0</ID>215 </input>
<input>
<ID>IN_1</ID>215 </input>
<output>
<ID>OUT</ID>211 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>388</ID>
<type>AA_TOGGLE</type>
<position>33.5,-200</position>
<output>
<ID>OUT_0</ID>206 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<wire>
<ID>193</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>40,-167.5,42.5,-167.5</points>
<connection>
<GID>362</GID>
<name>N_in0</name></connection>
<connection>
<GID>356</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>194</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>40,-174.5,42.5,-174.5</points>
<connection>
<GID>363</GID>
<name>N_in0</name></connection>
<intersection>40 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>40,-174.5,40,-174.5</points>
<connection>
<GID>357</GID>
<name>OUT</name></connection>
<intersection>-174.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>195</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>29.5,-166.5,34,-166.5</points>
<connection>
<GID>358</GID>
<name>OUT_0</name></connection>
<connection>
<GID>356</GID>
<name>IN_0</name></connection>
<intersection>33.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>33.5,-169.5,33.5,-166.5</points>
<connection>
<GID>454</GID>
<name>IN_0</name></connection>
<intersection>-166.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>25,-13,27.5,-13</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<connection>
<GID>4</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>25,-15,27.5,-15</points>
<connection>
<GID>2</GID>
<name>IN_1</name></connection>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>33.5,-14,36.5,-14</points>
<connection>
<GID>2</GID>
<name>OUT</name></connection>
<connection>
<GID>8</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>198</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>88.5,-166.5,93.5,-166.5</points>
<connection>
<GID>371</GID>
<name>IN_0</name></connection>
<intersection>88.5 7</intersection>
<intersection>90.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>90.5,-185.5,90.5,-166.5</points>
<intersection>-185.5 6</intersection>
<intersection>-180.5 4</intersection>
<intersection>-166.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>90.5,-180.5,100.5,-180.5</points>
<connection>
<GID>373</GID>
<name>IN_1</name></connection>
<intersection>90.5 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>90.5,-185.5,104.5,-185.5</points>
<connection>
<GID>374</GID>
<name>IN_1</name></connection>
<intersection>90.5 3</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>88.5,-166.5,88.5,-165.5</points>
<connection>
<GID>369</GID>
<name>OUT_0</name></connection>
<intersection>-166.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>54,-8,56.5,-8</points>
<connection>
<GID>26</GID>
<name>OUT_0</name></connection>
<connection>
<GID>24</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>199</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>108,-175.5,108,-173.5</points>
<intersection>-175.5 1</intersection>
<intersection>-173.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>108,-175.5,110,-175.5</points>
<connection>
<GID>375</GID>
<name>IN_0</name></connection>
<intersection>108 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>106.5,-173.5,108,-173.5</points>
<connection>
<GID>372</GID>
<name>OUT</name></connection>
<intersection>108 0</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>54,-10,56.5,-10</points>
<connection>
<GID>25</GID>
<name>OUT_0</name></connection>
<connection>
<GID>24</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>200</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>108,-179.5,108,-177.5</points>
<intersection>-179.5 1</intersection>
<intersection>-177.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>106.5,-179.5,108,-179.5</points>
<connection>
<GID>373</GID>
<name>OUT</name></connection>
<intersection>108 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>108,-177.5,110,-177.5</points>
<connection>
<GID>375</GID>
<name>IN_1</name></connection>
<intersection>108 0</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>54,-13.5,56.5,-13.5</points>
<connection>
<GID>22</GID>
<name>IN_0</name></connection>
<connection>
<GID>27</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>201</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>83,-183.5,83,-171</points>
<connection>
<GID>370</GID>
<name>OUT_0</name></connection>
<intersection>-183.5 3</intersection>
<intersection>-178.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>83,-178.5,100.5,-178.5</points>
<connection>
<GID>373</GID>
<name>IN_0</name></connection>
<intersection>83 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>83,-183.5,104.5,-183.5</points>
<connection>
<GID>374</GID>
<name>IN_0</name></connection>
<intersection>83 0</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>54,-15.5,56.5,-15.5</points>
<connection>
<GID>22</GID>
<name>IN_1</name></connection>
<connection>
<GID>28</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>202</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>93.5,-174.5,93.5,-170.5</points>
<connection>
<GID>371</GID>
<name>OUT_0</name></connection>
<intersection>-174.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>93.5,-174.5,100.5,-174.5</points>
<connection>
<GID>372</GID>
<name>IN_1</name></connection>
<intersection>93.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>25,-7.5,27.5,-7.5</points>
<connection>
<GID>10</GID>
<name>IN_0</name></connection>
<connection>
<GID>29</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>203</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>116,-176.5,120,-176.5</points>
<connection>
<GID>376</GID>
<name>N_in0</name></connection>
<connection>
<GID>375</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>25,-9.5,27.5,-9.5</points>
<connection>
<GID>10</GID>
<name>IN_1</name></connection>
<connection>
<GID>30</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>204</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>110.5,-184.5,114.5,-184.5</points>
<connection>
<GID>374</GID>
<name>OUT</name></connection>
<intersection>114.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>114.5,-186.5,114.5,-184.5</points>
<connection>
<GID>377</GID>
<name>N_in0</name></connection>
<intersection>-184.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>25,-3,27.5,-3</points>
<connection>
<GID>20</GID>
<name>IN_0</name></connection>
<connection>
<GID>31</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>205</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>78,-172.5,78,-166</points>
<connection>
<GID>368</GID>
<name>OUT_0</name></connection>
<intersection>-172.5 1</intersection>
<intersection>-167 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>78,-172.5,100.5,-172.5</points>
<connection>
<GID>372</GID>
<name>IN_0</name></connection>
<intersection>78 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>78,-167,83,-167</points>
<connection>
<GID>370</GID>
<name>IN_0</name></connection>
<intersection>78 0</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33.5,-3,33.5,-3</points>
<connection>
<GID>33</GID>
<name>N_in0</name></connection>
<connection>
<GID>20</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>206</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>33.5,-202,39.5,-202</points>
<connection>
<GID>388</GID>
<name>OUT_0</name></connection>
<connection>
<GID>389</GID>
<name>IN_1</name></connection>
<connection>
<GID>389</GID>
<name>IN_0</name></connection>
<intersection>35 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>35,-226,35,-202</points>
<intersection>-226 8</intersection>
<intersection>-218 6</intersection>
<intersection>-202 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>35,-218,48,-218</points>
<connection>
<GID>391</GID>
<name>IN_1</name></connection>
<intersection>35 5</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>35,-226,48.5,-226</points>
<connection>
<GID>392</GID>
<name>IN_1</name></connection>
<intersection>35 5</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33.5,-8.5,33.5,-8.5</points>
<connection>
<GID>35</GID>
<name>N_in0</name></connection>
<connection>
<GID>10</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>207</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56.5,-213.5,56.5,-212</points>
<intersection>-213.5 1</intersection>
<intersection>-212 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>56.5,-213.5,59.5,-213.5</points>
<connection>
<GID>394</GID>
<name>IN_0</name></connection>
<intersection>56.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>54,-212,56.5,-212</points>
<connection>
<GID>390</GID>
<name>OUT</name></connection>
<intersection>56.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>62.5,-9,64,-9</points>
<connection>
<GID>34</GID>
<name>N_in0</name></connection>
<connection>
<GID>24</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>208</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56.5,-217,56.5,-215.5</points>
<intersection>-217 1</intersection>
<intersection>-215.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>54,-217,56.5,-217</points>
<connection>
<GID>391</GID>
<name>OUT</name></connection>
<intersection>56.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>56.5,-215.5,59.5,-215.5</points>
<connection>
<GID>394</GID>
<name>IN_1</name></connection>
<intersection>56.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>209</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>54.5,-225,59.5,-225</points>
<connection>
<GID>392</GID>
<name>OUT</name></connection>
<intersection>59.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>59.5,-226,59.5,-224</points>
<connection>
<GID>393</GID>
<name>IN_1</name></connection>
<connection>
<GID>393</GID>
<name>IN_0</name></connection>
<intersection>-225 1</intersection></vsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>62.5,-14.5,64,-14.5</points>
<connection>
<GID>22</GID>
<name>OUT</name></connection>
<connection>
<GID>36</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19,-23.5,20.5,-23.5</points>
<connection>
<GID>55</GID>
<name>OUT_0</name></connection>
<intersection>20.5 10</intersection>
<intersection>20.5 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>20.5,-24.5,20.5,-22.5</points>
<connection>
<GID>53</GID>
<name>IN_1</name></connection>
<connection>
<GID>53</GID>
<name>IN_0</name></connection>
<intersection>-23.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>211</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29,-224,29,-209</points>
<connection>
<GID>387</GID>
<name>OUT</name></connection>
<intersection>-224 3</intersection>
<intersection>-216 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>29,-216,48,-216</points>
<connection>
<GID>391</GID>
<name>IN_0</name></connection>
<intersection>29 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>29,-224,48.5,-224</points>
<connection>
<GID>392</GID>
<name>IN_0</name></connection>
<intersection>29 0</intersection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26.5,-23.5,27.5,-23.5</points>
<connection>
<GID>53</GID>
<name>OUT</name></connection>
<connection>
<GID>57</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>212</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38.5,-213,38.5,-208</points>
<connection>
<GID>389</GID>
<name>OUT</name></connection>
<intersection>-213 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>38.5,-213,48,-213</points>
<connection>
<GID>390</GID>
<name>IN_1</name></connection>
<intersection>38.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>45,-25,45,-23</points>
<intersection>-25 3</intersection>
<intersection>-24 2</intersection>
<intersection>-23 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>45,-23,46.5,-23</points>
<connection>
<GID>61</GID>
<name>IN_0</name></connection>
<intersection>45 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>44,-24,45,-24</points>
<connection>
<GID>59</GID>
<name>OUT</name></connection>
<intersection>45 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>45,-25,46.5,-25</points>
<connection>
<GID>61</GID>
<name>IN_1</name></connection>
<intersection>45 0</intersection></hsegment></shape></wire>
<wire>
<ID>213</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>65.5,-214.5,68.5,-214.5</points>
<connection>
<GID>394</GID>
<name>OUT</name></connection>
<connection>
<GID>395</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38,-23,38,-23</points>
<connection>
<GID>62</GID>
<name>OUT_0</name></connection>
<connection>
<GID>59</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>214</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>65.5,-225,69,-225</points>
<connection>
<GID>393</GID>
<name>OUT</name></connection>
<connection>
<GID>396</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38,-25,38,-25</points>
<connection>
<GID>63</GID>
<name>OUT_0</name></connection>
<connection>
<GID>59</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>215</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>23.5,-211,23.5,-202</points>
<connection>
<GID>384</GID>
<name>OUT_0</name></connection>
<intersection>-211 1</intersection>
<intersection>-202.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>23.5,-211,48,-211</points>
<connection>
<GID>390</GID>
<name>IN_0</name></connection>
<intersection>23.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>23.5,-202.5,30,-202.5</points>
<intersection>23.5 0</intersection>
<intersection>28 4</intersection>
<intersection>30 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>30,-203,30,-202.5</points>
<connection>
<GID>387</GID>
<name>IN_0</name></connection>
<intersection>-202.5 2</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>28,-203,28,-202.5</points>
<connection>
<GID>387</GID>
<name>IN_1</name></connection>
<intersection>-202.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>52.5,-24,53.5,-24</points>
<connection>
<GID>64</GID>
<name>N_in0</name></connection>
<connection>
<GID>61</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>76.5,-25.5,76.5,-23.5</points>
<intersection>-25.5 1</intersection>
<intersection>-23.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>76.5,-25.5,78,-25.5</points>
<connection>
<GID>70</GID>
<name>IN_0</name></connection>
<intersection>76.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>75.5,-23.5,76.5,-23.5</points>
<connection>
<GID>66</GID>
<name>OUT</name></connection>
<intersection>76.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>217</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>98.5,-212.5,98.5,-202</points>
<connection>
<GID>409</GID>
<name>OUT_0</name></connection>
<intersection>-212.5 1</intersection>
<intersection>-204 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>98.5,-212.5,113,-212.5</points>
<connection>
<GID>404</GID>
<name>IN_1</name></connection>
<intersection>98.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>98.5,-204,103.5,-204</points>
<connection>
<GID>410</GID>
<name>IN_1</name></connection>
<connection>
<GID>410</GID>
<name>IN_0</name></connection>
<intersection>98.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>76.5,-29,76.5,-27.5</points>
<intersection>-29 2</intersection>
<intersection>-27.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>76.5,-27.5,78,-27.5</points>
<connection>
<GID>70</GID>
<name>IN_1</name></connection>
<intersection>76.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>75.5,-29,76.5,-29</points>
<connection>
<GID>68</GID>
<name>OUT</name></connection>
<intersection>76.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>218</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>102.5,-226.5,102.5,-210</points>
<connection>
<GID>410</GID>
<name>OUT</name></connection>
<intersection>-226.5 3</intersection>
<intersection>-217.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>102.5,-217.5,113,-217.5</points>
<connection>
<GID>405</GID>
<name>IN_1</name></connection>
<intersection>102.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>102.5,-226.5,112.5,-226.5</points>
<connection>
<GID>406</GID>
<name>IN_1</name></connection>
<intersection>102.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>219</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89,-224.5,89,-202</points>
<connection>
<GID>401</GID>
<name>OUT_0</name></connection>
<intersection>-224.5 6</intersection>
<intersection>-215.5 1</intersection>
<intersection>-204 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>89,-215.5,113,-215.5</points>
<connection>
<GID>405</GID>
<name>IN_0</name></connection>
<intersection>89 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>89,-204,94,-204</points>
<connection>
<GID>408</GID>
<name>IN_1</name></connection>
<connection>
<GID>408</GID>
<name>IN_0</name></connection>
<intersection>89 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>89,-224.5,112.5,-224.5</points>
<connection>
<GID>406</GID>
<name>IN_0</name></connection>
<intersection>89 0</intersection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>69,-24.5,69,-22.5</points>
<intersection>-24.5 1</intersection>
<intersection>-23.5 3</intersection>
<intersection>-22.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>69,-24.5,69.5,-24.5</points>
<connection>
<GID>66</GID>
<name>IN_1</name></connection>
<intersection>69 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>69,-22.5,69.5,-22.5</points>
<connection>
<GID>66</GID>
<name>IN_0</name></connection>
<intersection>69 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>67,-23.5,69,-23.5</points>
<connection>
<GID>71</GID>
<name>OUT_0</name></connection>
<intersection>69 0</intersection></hsegment></shape></wire>
<wire>
<ID>220</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>121,-213,121,-211.5</points>
<intersection>-213 2</intersection>
<intersection>-211.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>119,-211.5,121,-211.5</points>
<connection>
<GID>404</GID>
<name>OUT</name></connection>
<intersection>121 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>121,-213,123,-213</points>
<connection>
<GID>407</GID>
<name>IN_0</name></connection>
<intersection>121 0</intersection></hsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>69.5,-30,69.5,-28</points>
<connection>
<GID>68</GID>
<name>IN_1</name></connection>
<connection>
<GID>68</GID>
<name>IN_0</name></connection>
<intersection>-29 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>67,-29,69.5,-29</points>
<connection>
<GID>72</GID>
<name>OUT_0</name></connection>
<intersection>69.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>221</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>121,-216.5,121,-215</points>
<intersection>-216.5 1</intersection>
<intersection>-215 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>119,-216.5,121,-216.5</points>
<connection>
<GID>405</GID>
<name>OUT</name></connection>
<intersection>121 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>121,-215,123,-215</points>
<connection>
<GID>407</GID>
<name>IN_1</name></connection>
<intersection>121 0</intersection></hsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>84,-26.5,85,-26.5</points>
<connection>
<GID>70</GID>
<name>OUT</name></connection>
<connection>
<GID>74</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>222</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>118.5,-225.5,122.5,-225.5</points>
<connection>
<GID>412</GID>
<name>N_in0</name></connection>
<connection>
<GID>406</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>223</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>137.5,-214,140,-214</points>
<connection>
<GID>414</GID>
<name>OUT</name></connection>
<connection>
<GID>411</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>224</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>130,-215,130,-213</points>
<intersection>-215 3</intersection>
<intersection>-214 1</intersection>
<intersection>-213 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>129,-214,130,-214</points>
<connection>
<GID>407</GID>
<name>OUT</name></connection>
<intersection>130 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>130,-213,131.5,-213</points>
<connection>
<GID>414</GID>
<name>IN_0</name></connection>
<intersection>130 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>130,-215,131.5,-215</points>
<connection>
<GID>414</GID>
<name>IN_1</name></connection>
<intersection>130 0</intersection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37.5,-39,37.5,-36.5</points>
<intersection>-39 1</intersection>
<intersection>-36.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>37.5,-39,39,-39</points>
<connection>
<GID>79</GID>
<name>IN_0</name></connection>
<intersection>37.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>36.5,-36.5,37.5,-36.5</points>
<connection>
<GID>77</GID>
<name>OUT</name></connection>
<intersection>37.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>225</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>93,-211,93,-210</points>
<connection>
<GID>408</GID>
<name>OUT</name></connection>
<intersection>-211 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>93,-211,113,-211</points>
<intersection>93 0</intersection>
<intersection>113 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>113,-211,113,-210.5</points>
<connection>
<GID>404</GID>
<name>IN_0</name></connection>
<intersection>-211 1</intersection></vsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37.5,-43,37.5,-41</points>
<intersection>-43 1</intersection>
<intersection>-41 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>36,-43,37.5,-43</points>
<connection>
<GID>78</GID>
<name>OUT</name></connection>
<intersection>37.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>37.5,-41,39,-41</points>
<connection>
<GID>79</GID>
<name>IN_1</name></connection>
<intersection>37.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>226</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>53,-278.5,53,-274.5</points>
<intersection>-278.5 1</intersection>
<intersection>-274.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>53,-278.5,56,-278.5</points>
<connection>
<GID>426</GID>
<name>IN_0</name></connection>
<intersection>53 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>50,-274.5,53,-274.5</points>
<connection>
<GID>422</GID>
<name>OUT</name></connection>
<intersection>53 0</intersection></hsegment></shape></wire>
<wire>
<ID>227</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>50,-280.5,56,-280.5</points>
<connection>
<GID>423</GID>
<name>OUT</name></connection>
<connection>
<GID>426</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30,-42,30,-37.5</points>
<connection>
<GID>78</GID>
<name>IN_0</name></connection>
<intersection>-39.5 2</intersection>
<intersection>-37.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30,-37.5,30.5,-37.5</points>
<connection>
<GID>77</GID>
<name>IN_1</name></connection>
<intersection>30 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>28.5,-39.5,30,-39.5</points>
<connection>
<GID>76</GID>
<name>OUT</name></connection>
<intersection>30 0</intersection></hsegment></shape></wire>
<wire>
<ID>228</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>53,-286,53,-282.5</points>
<intersection>-286 1</intersection>
<intersection>-282.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50,-286,53,-286</points>
<connection>
<GID>424</GID>
<name>OUT</name></connection>
<intersection>53 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>53,-282.5,56,-282.5</points>
<connection>
<GID>426</GID>
<name>IN_2</name></connection>
<intersection>53 0</intersection></hsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22,-44,22,-40.5</points>
<intersection>-44 1</intersection>
<intersection>-42.5 2</intersection>
<intersection>-40.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>22,-44,30,-44</points>
<connection>
<GID>78</GID>
<name>IN_1</name></connection>
<intersection>22 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>20,-42.5,22,-42.5</points>
<connection>
<GID>85</GID>
<name>OUT_0</name></connection>
<intersection>22 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>22,-40.5,22.5,-40.5</points>
<connection>
<GID>76</GID>
<name>IN_1</name></connection>
<intersection>22 0</intersection></hsegment></shape></wire>
<wire>
<ID>229</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24.5,-285,24.5,-260</points>
<connection>
<GID>428</GID>
<name>OUT_0</name></connection>
<intersection>-285 5</intersection>
<intersection>-273.5 3</intersection>
<intersection>-261.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>24.5,-261.5,38,-261.5</points>
<connection>
<GID>420</GID>
<name>IN_0</name></connection>
<intersection>24.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>24.5,-273.5,44,-273.5</points>
<connection>
<GID>422</GID>
<name>IN_0</name></connection>
<intersection>24.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>24.5,-285,44,-285</points>
<connection>
<GID>424</GID>
<name>IN_0</name></connection>
<intersection>24.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>20,-35.5,30.5,-35.5</points>
<connection>
<GID>77</GID>
<name>IN_0</name></connection>
<connection>
<GID>73</GID>
<name>OUT_0</name></connection>
<intersection>21.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>21.5,-38.5,21.5,-35.5</points>
<intersection>-38.5 4</intersection>
<intersection>-35.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>21.5,-38.5,22.5,-38.5</points>
<connection>
<GID>76</GID>
<name>IN_0</name></connection>
<intersection>21.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>230</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28,-279.5,28,-260</points>
<connection>
<GID>429</GID>
<name>OUT_0</name></connection>
<intersection>-279.5 5</intersection>
<intersection>-275.5 3</intersection>
<intersection>-263.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>28,-263.5,38,-263.5</points>
<connection>
<GID>420</GID>
<name>IN_1</name></connection>
<intersection>28 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>28,-275.5,44,-275.5</points>
<connection>
<GID>422</GID>
<name>IN_1</name></connection>
<intersection>28 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>28,-279.5,44,-279.5</points>
<connection>
<GID>423</GID>
<name>IN_0</name></connection>
<intersection>28 0</intersection></hsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45,-40,47,-40</points>
<connection>
<GID>79</GID>
<name>OUT</name></connection>
<connection>
<GID>87</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>231</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31.5,-287,31.5,-260</points>
<connection>
<GID>430</GID>
<name>OUT_0</name></connection>
<intersection>-287 5</intersection>
<intersection>-281.5 3</intersection>
<intersection>-265.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>31.5,-265.5,38,-265.5</points>
<connection>
<GID>420</GID>
<name>IN_2</name></connection>
<intersection>31.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>31.5,-281.5,44,-281.5</points>
<connection>
<GID>423</GID>
<name>IN_1</name></connection>
<intersection>31.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>31.5,-287,44,-287</points>
<connection>
<GID>424</GID>
<name>IN_1</name></connection>
<intersection>31.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>91.5,-41.5,91.5,-37</points>
<intersection>-41.5 1</intersection>
<intersection>-37 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>91.5,-41.5,98.5,-41.5</points>
<connection>
<GID>83</GID>
<name>IN_0</name></connection>
<intersection>91.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>85,-37,91.5,-37</points>
<connection>
<GID>80</GID>
<name>OUT</name></connection>
<intersection>91.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>232</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>44,-263.5,49,-263.5</points>
<connection>
<GID>420</GID>
<name>OUT</name></connection>
<intersection>47 5</intersection>
<intersection>49 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>49,-263.5,49,-263</points>
<intersection>-263.5 1</intersection>
<intersection>-263 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>48,-263,49,-263</points>
<connection>
<GID>432</GID>
<name>N_in3</name></connection>
<intersection>49 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>47,-264,47,-263.5</points>
<connection>
<GID>432</GID>
<name>N_in0</name></connection>
<intersection>-263.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>96,-45.5,96,-43.5</points>
<intersection>-45.5 2</intersection>
<intersection>-43.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>96,-43.5,98.5,-43.5</points>
<connection>
<GID>83</GID>
<name>IN_1</name></connection>
<intersection>96 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>94.5,-45.5,96,-45.5</points>
<connection>
<GID>82</GID>
<name>OUT</name></connection>
<intersection>96 0</intersection></hsegment></shape></wire>
<wire>
<ID>233</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>62,-280.5,64.5,-280.5</points>
<connection>
<GID>433</GID>
<name>N_in0</name></connection>
<connection>
<GID>426</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>86.5,-44.5,86.5,-43</points>
<intersection>-44.5 1</intersection>
<intersection>-43 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>86.5,-44.5,88.5,-44.5</points>
<connection>
<GID>82</GID>
<name>IN_0</name></connection>
<intersection>86.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>85.5,-43,86.5,-43</points>
<connection>
<GID>81</GID>
<name>OUT</name></connection>
<intersection>86.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>234</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>33.5,-173.5,34,-173.5</points>
<connection>
<GID>454</GID>
<name>OUT_0</name></connection>
<connection>
<GID>357</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>86.5,-48,86.5,-46.5</points>
<intersection>-48 2</intersection>
<intersection>-46.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>86.5,-46.5,88.5,-46.5</points>
<connection>
<GID>82</GID>
<name>IN_1</name></connection>
<intersection>86.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>85,-48,86.5,-48</points>
<connection>
<GID>84</GID>
<name>OUT</name></connection>
<intersection>86.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>235</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>151.5,-278,151.5,-267</points>
<intersection>-278 1</intersection>
<intersection>-267 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>151.5,-278,160,-278</points>
<intersection>151.5 0</intersection>
<intersection>160 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>143,-267,151.5,-267</points>
<connection>
<GID>445</GID>
<name>OUT</name></connection>
<intersection>151.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>160,-279,160,-278</points>
<intersection>-279 4</intersection>
<intersection>-278 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>160,-279,162,-279</points>
<connection>
<GID>464</GID>
<name>IN_0</name></connection>
<intersection>160 3</intersection></hsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>77.5,-44,77.5,-36</points>
<intersection>-44 3</intersection>
<intersection>-42 2</intersection>
<intersection>-36 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>73.5,-36,79,-36</points>
<connection>
<GID>89</GID>
<name>OUT_0</name></connection>
<connection>
<GID>80</GID>
<name>IN_0</name></connection>
<intersection>77.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>77.5,-42,79.5,-42</points>
<connection>
<GID>81</GID>
<name>IN_0</name></connection>
<intersection>77.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>77.5,-44,79.5,-44</points>
<connection>
<GID>81</GID>
<name>IN_1</name></connection>
<intersection>77.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>236</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>150,-281,150,-275.5</points>
<intersection>-281 2</intersection>
<intersection>-275.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>144,-275.5,150,-275.5</points>
<connection>
<GID>446</GID>
<name>OUT</name></connection>
<intersection>150 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>150,-281,162,-281</points>
<connection>
<GID>464</GID>
<name>IN_1</name></connection>
<intersection>150 0</intersection></hsegment></shape></wire>
<wire>
<ID>237</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>150,-284,150,-283</points>
<intersection>-284 1</intersection>
<intersection>-283 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>143,-284,150,-284</points>
<intersection>143 3</intersection>
<intersection>150 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>150,-283,162,-283</points>
<connection>
<GID>464</GID>
<name>IN_2</name></connection>
<intersection>150 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>143,-284.5,143,-284</points>
<connection>
<GID>447</GID>
<name>OUT</name></connection>
<intersection>-284 1</intersection></vsegment></shape></wire>
<wire>
<ID>238</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>151.5,-294,151.5,-285</points>
<intersection>-294 1</intersection>
<intersection>-285 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>143,-294,151.5,-294</points>
<connection>
<GID>448</GID>
<name>OUT</name></connection>
<intersection>151.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>151.5,-285,162,-285</points>
<connection>
<GID>464</GID>
<name>IN_3</name></connection>
<intersection>151.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73.5,-38,79,-38</points>
<connection>
<GID>90</GID>
<name>OUT_0</name></connection>
<connection>
<GID>80</GID>
<name>IN_1</name></connection>
<intersection>78.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>78.5,-47,78.5,-38</points>
<intersection>-47 3</intersection>
<intersection>-38 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>78.5,-47,79,-47</points>
<connection>
<GID>84</GID>
<name>IN_0</name></connection>
<intersection>78.5 2</intersection>
<intersection>79 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>79,-49,79,-47</points>
<connection>
<GID>84</GID>
<name>IN_1</name></connection>
<intersection>-47 3</intersection></vsegment></shape></wire>
<wire>
<ID>239</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>156,-318.5,156,-308.5</points>
<intersection>-318.5 1</intersection>
<intersection>-308.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>156,-318.5,161,-318.5</points>
<connection>
<GID>465</GID>
<name>IN_0</name></connection>
<intersection>156 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>143,-308.5,156,-308.5</points>
<connection>
<GID>449</GID>
<name>OUT</name></connection>
<intersection>156 0</intersection></hsegment></shape></wire>
<wire>
<ID>46</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>104.5,-42.5,105.5,-42.5</points>
<connection>
<GID>83</GID>
<name>OUT</name></connection>
<connection>
<GID>97</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>240</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>152,-320.5,152,-318</points>
<intersection>-320.5 2</intersection>
<intersection>-318 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>143,-318,152,-318</points>
<connection>
<GID>450</GID>
<name>OUT</name></connection>
<intersection>152 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>152,-320.5,161,-320.5</points>
<connection>
<GID>465</GID>
<name>IN_1</name></connection>
<intersection>152 0</intersection></hsegment></shape></wire>
<wire>
<ID>241</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>152,-327,152,-322.5</points>
<intersection>-327 1</intersection>
<intersection>-322.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>143,-327,152,-327</points>
<connection>
<GID>451</GID>
<name>OUT</name></connection>
<intersection>152 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>152,-322.5,161,-322.5</points>
<connection>
<GID>465</GID>
<name>IN_2</name></connection>
<intersection>152 0</intersection></hsegment></shape></wire>
<wire>
<ID>242</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>156.5,-336.5,156.5,-324.5</points>
<intersection>-336.5 1</intersection>
<intersection>-324.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>143,-336.5,156.5,-336.5</points>
<connection>
<GID>452</GID>
<name>OUT</name></connection>
<intersection>156.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>156.5,-324.5,161,-324.5</points>
<connection>
<GID>465</GID>
<name>IN_3</name></connection>
<intersection>156.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>50</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>86.5,-8.5,89,-8.5</points>
<connection>
<GID>102</GID>
<name>OUT_0</name></connection>
<connection>
<GID>110</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>244</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>111,-327,111,-253</points>
<connection>
<GID>457</GID>
<name>OUT_0</name></connection>
<intersection>-327 10</intersection>
<intersection>-318 8</intersection>
<intersection>-294 6</intersection>
<intersection>-275.5 3</intersection>
<intersection>-255 4</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>111,-275.5,138,-275.5</points>
<connection>
<GID>446</GID>
<name>IN_1</name></connection>
<intersection>111 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>111,-255,116,-255</points>
<connection>
<GID>461</GID>
<name>IN_0</name></connection>
<intersection>111 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>111,-294,137,-294</points>
<connection>
<GID>448</GID>
<name>IN_1</name></connection>
<intersection>111 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>111,-318,137,-318</points>
<connection>
<GID>450</GID>
<name>IN_1</name></connection>
<intersection>111 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>111,-327,137,-327</points>
<connection>
<GID>451</GID>
<name>IN_1</name></connection>
<intersection>111 0</intersection></hsegment></shape></wire>
<wire>
<ID>51</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>86.5,-10.5,89,-10.5</points>
<connection>
<GID>101</GID>
<name>OUT_0</name></connection>
<connection>
<GID>110</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>52</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>95,-9.5,96.5,-9.5</points>
<connection>
<GID>103</GID>
<name>N_in0</name></connection>
<connection>
<GID>110</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>246</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>103,-316,103,-259</points>
<connection>
<GID>460</GID>
<name>OUT_0</name></connection>
<intersection>-316 5</intersection>
<intersection>-273.5 3</intersection>
<intersection>-265 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>103,-265,137,-265</points>
<connection>
<GID>445</GID>
<name>IN_0</name></connection>
<intersection>103 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>103,-273.5,138,-273.5</points>
<connection>
<GID>446</GID>
<name>IN_0</name></connection>
<intersection>103 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>103,-316,137,-316</points>
<connection>
<GID>450</GID>
<name>IN_0</name></connection>
<intersection>103 0</intersection></hsegment></shape></wire>
<wire>
<ID>247</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>116,-308.5,116,-259</points>
<connection>
<GID>461</GID>
<name>OUT_0</name></connection>
<intersection>-308.5 5</intersection>
<intersection>-284.5 3</intersection>
<intersection>-267 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>116,-267,137,-267</points>
<connection>
<GID>445</GID>
<name>IN_1</name></connection>
<intersection>116 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>116,-284.5,137,-284.5</points>
<connection>
<GID>447</GID>
<name>IN_1</name></connection>
<intersection>116 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>116,-308.5,137,-308.5</points>
<connection>
<GID>449</GID>
<name>IN_1</name></connection>
<intersection>116 0</intersection></hsegment></shape></wire>
<wire>
<ID>248</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>122.5,-320,122.5,-253</points>
<connection>
<GID>458</GID>
<name>OUT_0</name></connection>
<intersection>-320 8</intersection>
<intersection>-310.5 6</intersection>
<intersection>-296 4</intersection>
<intersection>-269 1</intersection>
<intersection>-255 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>122.5,-269,137,-269</points>
<connection>
<GID>445</GID>
<name>IN_2</name></connection>
<intersection>122.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>122.5,-255,128,-255</points>
<connection>
<GID>462</GID>
<name>IN_0</name></connection>
<intersection>122.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>122.5,-296,137,-296</points>
<connection>
<GID>448</GID>
<name>IN_2</name></connection>
<intersection>122.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>122.5,-310.5,137,-310.5</points>
<connection>
<GID>449</GID>
<name>IN_2</name></connection>
<intersection>122.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>122.5,-320,137,-320</points>
<connection>
<GID>450</GID>
<name>IN_2</name></connection>
<intersection>122.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>249</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>128,-329,128,-259</points>
<connection>
<GID>462</GID>
<name>OUT_0</name></connection>
<intersection>-329 5</intersection>
<intersection>-286.5 3</intersection>
<intersection>-277.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>128,-277.5,138,-277.5</points>
<connection>
<GID>446</GID>
<name>IN_2</name></connection>
<intersection>128 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>128,-286.5,137,-286.5</points>
<connection>
<GID>447</GID>
<name>IN_2</name></connection>
<intersection>128 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>128,-329,137,-329</points>
<connection>
<GID>451</GID>
<name>IN_2</name></connection>
<intersection>128 0</intersection></hsegment></shape></wire>
<wire>
<ID>56</ID>
<shape>
<hsegment>
<ID>4</ID>
<points>86.5,-14,89.5,-14</points>
<connection>
<GID>112</GID>
<name>IN_0</name></connection>
<intersection>86.5 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>86.5,-14,86.5,-13.5</points>
<connection>
<GID>114</GID>
<name>OUT_0</name></connection>
<intersection>-14 4</intersection></vsegment></shape></wire>
<wire>
<ID>250</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>99,-325,99,-253</points>
<connection>
<GID>456</GID>
<name>OUT_0</name></connection>
<intersection>-325 8</intersection>
<intersection>-306.5 6</intersection>
<intersection>-292 4</intersection>
<intersection>-282.5 1</intersection>
<intersection>-255 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>99,-282.5,137,-282.5</points>
<connection>
<GID>447</GID>
<name>IN_0</name></connection>
<intersection>99 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>99,-255,103,-255</points>
<connection>
<GID>460</GID>
<name>IN_0</name></connection>
<intersection>99 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>99,-292,137,-292</points>
<connection>
<GID>448</GID>
<name>IN_0</name></connection>
<intersection>99 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>99,-306.5,137,-306.5</points>
<connection>
<GID>449</GID>
<name>IN_0</name></connection>
<intersection>99 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>99,-325,137,-325</points>
<connection>
<GID>451</GID>
<name>IN_0</name></connection>
<intersection>99 0</intersection></hsegment></shape></wire>
<wire>
<ID>63</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>86.5,-16,89.5,-16</points>
<connection>
<GID>113</GID>
<name>OUT_0</name></connection>
<connection>
<GID>112</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>65</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>95.5,-15,97,-15</points>
<connection>
<GID>115</GID>
<name>N_in0</name></connection>
<connection>
<GID>112</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>79</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32.5,-77,32.5,-73</points>
<intersection>-77 6</intersection>
<intersection>-75 4</intersection>
<intersection>-73 5</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>31.5,-75,32.5,-75</points>
<connection>
<GID>180</GID>
<name>OUT</name></connection>
<intersection>32.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>32.5,-73,35,-73</points>
<connection>
<GID>181</GID>
<name>IN_1</name></connection>
<intersection>32.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>32.5,-77,34.5,-77</points>
<connection>
<GID>182</GID>
<name>IN_0</name></connection>
<intersection>32.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>80</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>22.5,-79,34.5,-79</points>
<connection>
<GID>182</GID>
<name>IN_1</name></connection>
<connection>
<GID>159</GID>
<name>OUT_0</name></connection>
<intersection>25.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>25.5,-79,25.5,-76</points>
<connection>
<GID>180</GID>
<name>IN_1</name></connection>
<intersection>-79 2</intersection></vsegment></shape></wire>
<wire>
<ID>81</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>22.5,-71,35,-71</points>
<connection>
<GID>148</GID>
<name>OUT_0</name></connection>
<connection>
<GID>181</GID>
<name>IN_0</name></connection>
<intersection>25.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>25.5,-74,25.5,-71</points>
<connection>
<GID>180</GID>
<name>IN_0</name></connection>
<intersection>-71 1</intersection></vsegment></shape></wire>
<wire>
<ID>90</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22,-60,22,-58</points>
<intersection>-60 3</intersection>
<intersection>-59 2</intersection>
<intersection>-58 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>22,-58,23,-58</points>
<connection>
<GID>174</GID>
<name>IN_0</name></connection>
<intersection>22 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>21.5,-59,22,-59</points>
<connection>
<GID>136</GID>
<name>OUT_0</name></connection>
<intersection>22 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>22,-60,23,-60</points>
<connection>
<GID>174</GID>
<name>IN_1</name></connection>
<intersection>22 0</intersection></hsegment></shape></wire>
<wire>
<ID>91</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>29,-59,30,-59</points>
<connection>
<GID>137</GID>
<name>N_in0</name></connection>
<connection>
<GID>174</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>92</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>48.5,-60.5,48.5,-58.5</points>
<intersection>-60.5 3</intersection>
<intersection>-59.5 1</intersection>
<intersection>-58.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>48,-59.5,48.5,-59.5</points>
<connection>
<GID>175</GID>
<name>OUT</name></connection>
<intersection>48.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>48.5,-58.5,49,-58.5</points>
<connection>
<GID>176</GID>
<name>IN_0</name></connection>
<intersection>48.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>48.5,-60.5,49,-60.5</points>
<connection>
<GID>176</GID>
<name>IN_1</name></connection>
<intersection>48.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>93</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>55,-59.5,56,-59.5</points>
<connection>
<GID>142</GID>
<name>N_in0</name></connection>
<connection>
<GID>176</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>94</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>40.5,-58.5,42,-58.5</points>
<connection>
<GID>140</GID>
<name>OUT_0</name></connection>
<connection>
<GID>175</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>95</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>40.5,-60.5,42,-60.5</points>
<connection>
<GID>141</GID>
<name>OUT_0</name></connection>
<connection>
<GID>175</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>96</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>71.5,-59.5,71.5,-57.5</points>
<intersection>-59.5 3</intersection>
<intersection>-59 1</intersection>
<intersection>-57.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>69.5,-59,71.5,-59</points>
<connection>
<GID>146</GID>
<name>OUT_0</name></connection>
<intersection>71.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71.5,-57.5,72,-57.5</points>
<connection>
<GID>177</GID>
<name>IN_0</name></connection>
<intersection>71.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>71.5,-59.5,72,-59.5</points>
<connection>
<GID>177</GID>
<name>IN_1</name></connection>
<intersection>71.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>97</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>70.5,-65.5,70.5,-63.5</points>
<intersection>-65.5 3</intersection>
<intersection>-64.5 2</intersection>
<intersection>-63.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>70.5,-63.5,72,-63.5</points>
<connection>
<GID>178</GID>
<name>IN_0</name></connection>
<intersection>70.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>69.5,-64.5,70.5,-64.5</points>
<connection>
<GID>147</GID>
<name>OUT_0</name></connection>
<intersection>70.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>70.5,-65.5,72,-65.5</points>
<connection>
<GID>178</GID>
<name>IN_1</name></connection>
<intersection>70.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>98</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>79,-61,79,-58.5</points>
<intersection>-61 1</intersection>
<intersection>-58.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>79,-61,80.5,-61</points>
<connection>
<GID>179</GID>
<name>IN_0</name></connection>
<intersection>79 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>78,-58.5,79,-58.5</points>
<connection>
<GID>177</GID>
<name>OUT</name></connection>
<intersection>79 0</intersection></hsegment></shape></wire>
<wire>
<ID>99</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>79,-64.5,79,-63</points>
<intersection>-64.5 1</intersection>
<intersection>-63 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>78,-64.5,79,-64.5</points>
<connection>
<GID>178</GID>
<name>OUT</name></connection>
<intersection>79 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>79,-63,80.5,-63</points>
<connection>
<GID>179</GID>
<name>IN_1</name></connection>
<intersection>79 0</intersection></hsegment></shape></wire>
<wire>
<ID>100</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>86.5,-62,87.5,-62</points>
<connection>
<GID>149</GID>
<name>N_in0</name></connection>
<connection>
<GID>179</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>101</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>41.5,-74.5,41.5,-72</points>
<intersection>-74.5 1</intersection>
<intersection>-72 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>41.5,-74.5,42.5,-74.5</points>
<connection>
<GID>183</GID>
<name>IN_0</name></connection>
<intersection>41.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>41,-72,41.5,-72</points>
<connection>
<GID>181</GID>
<name>OUT</name></connection>
<intersection>41.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>102</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>41.5,-78,41.5,-76.5</points>
<intersection>-78 1</intersection>
<intersection>-76.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>40.5,-78,41.5,-78</points>
<connection>
<GID>182</GID>
<name>OUT</name></connection>
<intersection>41.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>41.5,-76.5,42.5,-76.5</points>
<connection>
<GID>183</GID>
<name>IN_1</name></connection>
<intersection>41.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>103</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>48.5,-75.5,49.5,-75.5</points>
<connection>
<GID>160</GID>
<name>N_in0</name></connection>
<connection>
<GID>183</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>110</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>75.5,-78.5,75.5,-74.5</points>
<intersection>-78.5 6</intersection>
<intersection>-76.5 4</intersection>
<intersection>-74.5 5</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>74.5,-76.5,75.5,-76.5</points>
<connection>
<GID>198</GID>
<name>OUT</name></connection>
<intersection>75.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>75.5,-74.5,78,-74.5</points>
<connection>
<GID>199</GID>
<name>IN_1</name></connection>
<intersection>75.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>75.5,-78.5,77.5,-78.5</points>
<connection>
<GID>200</GID>
<name>IN_0</name></connection>
<intersection>75.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>111</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>65.5,-80.5,77.5,-80.5</points>
<connection>
<GID>194</GID>
<name>OUT_0</name></connection>
<connection>
<GID>200</GID>
<name>IN_1</name></connection>
<intersection>68.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>68.5,-80.5,68.5,-77.5</points>
<connection>
<GID>198</GID>
<name>IN_1</name></connection>
<intersection>-80.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>112</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>65.5,-72.5,78,-72.5</points>
<connection>
<GID>193</GID>
<name>OUT_0</name></connection>
<connection>
<GID>199</GID>
<name>IN_0</name></connection>
<intersection>68.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>68.5,-75.5,68.5,-72.5</points>
<connection>
<GID>198</GID>
<name>IN_0</name></connection>
<intersection>-72.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>113</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>84.5,-76,84.5,-73.5</points>
<intersection>-76 1</intersection>
<intersection>-73.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>84.5,-76,85.5,-76</points>
<connection>
<GID>201</GID>
<name>IN_0</name></connection>
<intersection>84.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>84,-73.5,84.5,-73.5</points>
<connection>
<GID>199</GID>
<name>OUT</name></connection>
<intersection>84.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>114</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>84.5,-79.5,84.5,-78</points>
<intersection>-79.5 1</intersection>
<intersection>-78 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>83.5,-79.5,84.5,-79.5</points>
<connection>
<GID>200</GID>
<name>OUT</name></connection>
<intersection>84.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>84.5,-78,85.5,-78</points>
<connection>
<GID>201</GID>
<name>IN_1</name></connection>
<intersection>84.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>116</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>92.5,-78,92.5,-76</points>
<intersection>-78 3</intersection>
<intersection>-77 1</intersection>
<intersection>-76 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>91.5,-77,92.5,-77</points>
<connection>
<GID>201</GID>
<name>OUT</name></connection>
<intersection>92.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>92.5,-76,93.5,-76</points>
<connection>
<GID>202</GID>
<name>IN_0</name></connection>
<intersection>92.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>92.5,-78,93.5,-78</points>
<connection>
<GID>202</GID>
<name>IN_1</name></connection>
<intersection>92.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>117</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>99.5,-77,101,-77</points>
<connection>
<GID>195</GID>
<name>N_in0</name></connection>
<connection>
<GID>202</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>118</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>23.5,-95.5,28,-95.5</points>
<connection>
<GID>215</GID>
<name>IN_0</name></connection>
<connection>
<GID>218</GID>
<name>OUT_0</name></connection>
<intersection>26.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>26.5,-102.5,26.5,-95.5</points>
<intersection>-102.5 5</intersection>
<intersection>-95.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>26.5,-102.5,28,-102.5</points>
<connection>
<GID>217</GID>
<name>IN_0</name></connection>
<intersection>26.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>119</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25,-104.5,25,-97.5</points>
<intersection>-104.5 3</intersection>
<intersection>-98.5 1</intersection>
<intersection>-97.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>23.5,-98.5,25,-98.5</points>
<connection>
<GID>220</GID>
<name>OUT_0</name></connection>
<intersection>25 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>25,-97.5,28,-97.5</points>
<connection>
<GID>215</GID>
<name>IN_1</name></connection>
<intersection>25 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>25,-104.5,28,-104.5</points>
<connection>
<GID>217</GID>
<name>IN_1</name></connection>
<intersection>25 0</intersection></hsegment></shape></wire>
<wire>
<ID>120</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>34,-96.5,36.5,-96.5</points>
<connection>
<GID>215</GID>
<name>OUT</name></connection>
<connection>
<GID>223</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>122</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>34,-103.5,36.5,-103.5</points>
<connection>
<GID>225</GID>
<name>N_in0</name></connection>
<connection>
<GID>217</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>123</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>66,-111,66,-94</points>
<intersection>-111 13</intersection>
<intersection>-100 3</intersection>
<intersection>-94 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>63.5,-94,68.5,-94</points>
<intersection>63.5 11</intersection>
<intersection>66 0</intersection>
<intersection>68.5 14</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>66,-100,86,-100</points>
<connection>
<GID>234</GID>
<name>IN_0</name></connection>
<intersection>66 0</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>63.5,-94,63.5,-93.5</points>
<connection>
<GID>227</GID>
<name>OUT_0</name></connection>
<intersection>-94 2</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>66,-111,90,-111</points>
<connection>
<GID>236</GID>
<name>IN_0</name></connection>
<intersection>66 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>68.5,-94.5,68.5,-94</points>
<connection>
<GID>230</GID>
<name>IN_0</name></connection>
<intersection>-94 2</intersection></vsegment></shape></wire>
<wire>
<ID>124</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>74,-94,79,-94</points>
<connection>
<GID>232</GID>
<name>IN_0</name></connection>
<intersection>74 7</intersection>
<intersection>76 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>76,-113,76,-94</points>
<intersection>-113 6</intersection>
<intersection>-108 4</intersection>
<intersection>-94 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>76,-108,86,-108</points>
<connection>
<GID>235</GID>
<name>IN_1</name></connection>
<intersection>76 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>76,-113,90,-113</points>
<connection>
<GID>236</GID>
<name>IN_1</name></connection>
<intersection>76 3</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>74,-94,74,-93</points>
<connection>
<GID>228</GID>
<name>OUT_0</name></connection>
<intersection>-94 1</intersection></vsegment></shape></wire>
<wire>
<ID>125</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>93.5,-103,93.5,-101</points>
<intersection>-103 1</intersection>
<intersection>-101 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>93.5,-103,95.5,-103</points>
<connection>
<GID>238</GID>
<name>IN_0</name></connection>
<intersection>93.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>92,-101,93.5,-101</points>
<connection>
<GID>234</GID>
<name>OUT</name></connection>
<intersection>93.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>126</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>93.5,-107,93.5,-105</points>
<intersection>-107 1</intersection>
<intersection>-105 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>92,-107,93.5,-107</points>
<connection>
<GID>235</GID>
<name>OUT</name></connection>
<intersection>93.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>93.5,-105,95.5,-105</points>
<connection>
<GID>238</GID>
<name>IN_1</name></connection>
<intersection>93.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>127</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>68.5,-106,68.5,-98.5</points>
<connection>
<GID>230</GID>
<name>OUT_0</name></connection>
<intersection>-106 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>68.5,-106,86,-106</points>
<connection>
<GID>235</GID>
<name>IN_0</name></connection>
<intersection>68.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>128</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>79,-102,79,-98</points>
<connection>
<GID>232</GID>
<name>OUT_0</name></connection>
<intersection>-102 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>79,-102,86,-102</points>
<connection>
<GID>234</GID>
<name>IN_1</name></connection>
<intersection>79 0</intersection></hsegment></shape></wire>
<wire>
<ID>129</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>101.5,-104,105.5,-104</points>
<connection>
<GID>240</GID>
<name>N_in0</name></connection>
<connection>
<GID>238</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>130</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>96,-112,100,-112</points>
<connection>
<GID>236</GID>
<name>OUT</name></connection>
<intersection>100 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>100,-114,100,-112</points>
<connection>
<GID>242</GID>
<name>N_in0</name></connection>
<intersection>-112 1</intersection></vsegment></shape></wire>
<wire>
<ID>152</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>27.5,-124,33.5,-124</points>
<connection>
<GID>301</GID>
<name>IN_1</name></connection>
<connection>
<GID>301</GID>
<name>IN_0</name></connection>
<connection>
<GID>300</GID>
<name>OUT_0</name></connection>
<intersection>29 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>29,-148,29,-124</points>
<intersection>-148 8</intersection>
<intersection>-140 6</intersection>
<intersection>-124 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>29,-140,42,-140</points>
<connection>
<GID>303</GID>
<name>IN_1</name></connection>
<intersection>29 5</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>29,-148,42.5,-148</points>
<connection>
<GID>304</GID>
<name>IN_1</name></connection>
<intersection>29 5</intersection></hsegment></shape></wire>
<wire>
<ID>153</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50.5,-135.5,50.5,-134</points>
<intersection>-135.5 1</intersection>
<intersection>-134 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50.5,-135.5,53.5,-135.5</points>
<connection>
<GID>306</GID>
<name>IN_0</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>48,-134,50.5,-134</points>
<connection>
<GID>302</GID>
<name>OUT</name></connection>
<intersection>50.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>154</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50.5,-139,50.5,-137.5</points>
<intersection>-139 1</intersection>
<intersection>-137.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>48,-139,50.5,-139</points>
<connection>
<GID>303</GID>
<name>OUT</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>50.5,-137.5,53.5,-137.5</points>
<connection>
<GID>306</GID>
<name>IN_1</name></connection>
<intersection>50.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>155</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>48.5,-147,53.5,-147</points>
<connection>
<GID>304</GID>
<name>OUT</name></connection>
<intersection>53.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>53.5,-148,53.5,-146</points>
<connection>
<GID>305</GID>
<name>IN_1</name></connection>
<connection>
<GID>305</GID>
<name>IN_0</name></connection>
<intersection>-147 1</intersection></vsegment></shape></wire>
<wire>
<ID>156</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>17.5,-124,24,-124</points>
<connection>
<GID>296</GID>
<name>OUT_0</name></connection>
<intersection>19 3</intersection>
<intersection>22 4</intersection>
<intersection>24 7</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>19,-146,19,-124</points>
<intersection>-146 9</intersection>
<intersection>-133 5</intersection>
<intersection>-124 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>22,-124.5,22,-124</points>
<connection>
<GID>299</GID>
<name>IN_1</name></connection>
<intersection>-124 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>19,-133,42,-133</points>
<connection>
<GID>302</GID>
<name>IN_0</name></connection>
<intersection>19 3</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>24,-124.5,24,-124</points>
<connection>
<GID>299</GID>
<name>IN_0</name></connection>
<intersection>-124 1</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>19,-146,42.5,-146</points>
<connection>
<GID>304</GID>
<name>IN_0</name></connection>
<intersection>19 3</intersection></hsegment></shape></wire>
<wire>
<ID>157</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>23,-138,23,-130.5</points>
<connection>
<GID>299</GID>
<name>OUT</name></connection>
<intersection>-138 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>23,-138,42,-138</points>
<connection>
<GID>303</GID>
<name>IN_0</name></connection>
<intersection>23 0</intersection></hsegment></shape></wire>
<wire>
<ID>158</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32.5,-135,32.5,-130</points>
<connection>
<GID>301</GID>
<name>OUT</name></connection>
<intersection>-135 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>32.5,-135,42,-135</points>
<connection>
<GID>302</GID>
<name>IN_1</name></connection>
<intersection>32.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>159</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>59.5,-136.5,62.5,-136.5</points>
<connection>
<GID>307</GID>
<name>N_in0</name></connection>
<connection>
<GID>306</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>160</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>59.5,-147,63,-147</points>
<connection>
<GID>308</GID>
<name>N_in0</name></connection>
<connection>
<GID>305</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>181</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>81.5,-149,81.5,-134.5</points>
<connection>
<GID>347</GID>
<name>OUT</name></connection>
<intersection>-149 3</intersection>
<intersection>-135 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>81.5,-135,101.5,-135</points>
<connection>
<GID>327</GID>
<name>IN_0</name></connection>
<intersection>81.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>81.5,-149,101,-149</points>
<connection>
<GID>344</GID>
<name>IN_0</name></connection>
<intersection>81.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>183</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>87,-137,87,-126.5</points>
<connection>
<GID>348</GID>
<name>OUT_0</name></connection>
<intersection>-137 1</intersection>
<intersection>-128.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>87,-137,101.5,-137</points>
<connection>
<GID>327</GID>
<name>IN_1</name></connection>
<intersection>87 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>87,-128.5,92,-128.5</points>
<connection>
<GID>349</GID>
<name>IN_1</name></connection>
<connection>
<GID>349</GID>
<name>IN_0</name></connection>
<intersection>87 0</intersection></hsegment></shape></wire>
<wire>
<ID>184</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>91,-151,91,-134.5</points>
<connection>
<GID>349</GID>
<name>OUT</name></connection>
<intersection>-151 3</intersection>
<intersection>-142 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>91,-142,101.5,-142</points>
<connection>
<GID>343</GID>
<name>IN_1</name></connection>
<intersection>91 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>91,-151,101,-151</points>
<connection>
<GID>344</GID>
<name>IN_1</name></connection>
<intersection>91 0</intersection></hsegment></shape></wire>
<wire>
<ID>185</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>77,-140,77,-126.5</points>
<connection>
<GID>311</GID>
<name>OUT_0</name></connection>
<intersection>-140 1</intersection>
<intersection>-128.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>77,-140,101.5,-140</points>
<connection>
<GID>343</GID>
<name>IN_0</name></connection>
<intersection>77 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>77,-128.5,82.5,-128.5</points>
<connection>
<GID>347</GID>
<name>IN_0</name></connection>
<connection>
<GID>347</GID>
<name>IN_1</name></connection>
<intersection>77 0</intersection></hsegment></shape></wire>
<wire>
<ID>186</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>109.5,-137.5,109.5,-136</points>
<intersection>-137.5 2</intersection>
<intersection>-136 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>107.5,-136,109.5,-136</points>
<connection>
<GID>327</GID>
<name>OUT</name></connection>
<intersection>109.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>109.5,-137.5,111.5,-137.5</points>
<connection>
<GID>345</GID>
<name>IN_0</name></connection>
<intersection>109.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>187</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>109.5,-141,109.5,-139.5</points>
<intersection>-141 1</intersection>
<intersection>-139.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>107.5,-141,109.5,-141</points>
<connection>
<GID>343</GID>
<name>OUT</name></connection>
<intersection>109.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>109.5,-139.5,111.5,-139.5</points>
<connection>
<GID>345</GID>
<name>IN_1</name></connection>
<intersection>109.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>188</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>107,-150,111,-150</points>
<connection>
<GID>344</GID>
<name>OUT</name></connection>
<connection>
<GID>351</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>189</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>126,-138.5,128.5,-138.5</points>
<connection>
<GID>350</GID>
<name>N_in0</name></connection>
<connection>
<GID>353</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>190</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>118.5,-139.5,118.5,-137.5</points>
<intersection>-139.5 3</intersection>
<intersection>-138.5 1</intersection>
<intersection>-137.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>117.5,-138.5,118.5,-138.5</points>
<connection>
<GID>345</GID>
<name>OUT</name></connection>
<intersection>118.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>118.5,-137.5,120,-137.5</points>
<connection>
<GID>353</GID>
<name>IN_0</name></connection>
<intersection>118.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>118.5,-139.5,120,-139.5</points>
<connection>
<GID>353</GID>
<name>IN_1</name></connection>
<intersection>118.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>192</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31,-175.5,31,-168.5</points>
<intersection>-175.5 3</intersection>
<intersection>-169.5 1</intersection>
<intersection>-168.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>29.5,-169.5,31,-169.5</points>
<connection>
<GID>360</GID>
<name>OUT_0</name></connection>
<intersection>31 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>31,-168.5,34,-168.5</points>
<connection>
<GID>356</GID>
<name>IN_1</name></connection>
<intersection>31 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>31,-175.5,34,-175.5</points>
<connection>
<GID>357</GID>
<name>IN_1</name></connection>
<intersection>31 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,0,145.8,-73.7</PageViewport></page 1>
<page 2>
<PageViewport>0,0,145.8,-73.7</PageViewport></page 2>
<page 3>
<PageViewport>0,0,145.8,-73.7</PageViewport></page 3>
<page 4>
<PageViewport>0,0,145.8,-73.7</PageViewport></page 4>
<page 5>
<PageViewport>0,0,145.8,-73.7</PageViewport></page 5>
<page 6>
<PageViewport>0,0,145.8,-73.7</PageViewport></page 6>
<page 7>
<PageViewport>0,0,145.8,-73.7</PageViewport></page 7>
<page 8>
<PageViewport>0,0,145.8,-73.7</PageViewport></page 8>
<page 9>
<PageViewport>0,0,145.8,-73.7</PageViewport></page 9></circuit>