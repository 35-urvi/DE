<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-91.3284,76.9034,297.472,-119.63</PageViewport>
<gate>
<ID>193</ID>
<type>AA_AND3</type>
<position>64,-71.5</position>
<input>
<ID>IN_0</ID>80 </input>
<input>
<ID>IN_1</ID>83 </input>
<input>
<ID>IN_2</ID>79 </input>
<output>
<ID>OUT</ID>87 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>194</ID>
<type>AA_AND3</type>
<position>64,-79.5</position>
<input>
<ID>IN_0</ID>81 </input>
<input>
<ID>IN_1</ID>82 </input>
<input>
<ID>IN_2</ID>79 </input>
<output>
<ID>OUT</ID>84 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>195</ID>
<type>AA_AND3</type>
<position>64,-87.5</position>
<input>
<ID>IN_0</ID>81 </input>
<input>
<ID>IN_1</ID>83 </input>
<input>
<ID>IN_2</ID>79 </input>
<output>
<ID>OUT</ID>85 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>2</ID>
<type>AA_MUX_2x1</type>
<position>24,-8</position>
<input>
<ID>IN_0</ID>2 </input>
<input>
<ID>IN_1</ID>1 </input>
<output>
<ID>OUT</ID>3 </output>
<input>
<ID>SEL_0</ID>4 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>196</ID>
<type>AA_LABEL</type>
<position>35.5,-50</position>
<gparam>LABEL_TEXT S0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>197</ID>
<type>AA_LABEL</type>
<position>26,-50</position>
<gparam>LABEL_TEXT S1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>4</ID>
<type>AA_TOGGLE</type>
<position>17.5,-7</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>198</ID>
<type>AA_LABEL</type>
<position>43.5,-50</position>
<gparam>LABEL_TEXT Din</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>199</ID>
<type>GA_LED</type>
<position>76.5,-63.5</position>
<input>
<ID>N_in0</ID>86 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>6</ID>
<type>AA_TOGGLE</type>
<position>20,-9</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>200</ID>
<type>GA_LED</type>
<position>76.5,-71.5</position>
<input>
<ID>N_in0</ID>87 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>201</ID>
<type>GA_LED</type>
<position>77,-79.5</position>
<input>
<ID>N_in0</ID>84 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>8</ID>
<type>GA_LED</type>
<position>27,-8</position>
<input>
<ID>N_in0</ID>3 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>202</ID>
<type>GA_LED</type>
<position>77,-87.5</position>
<input>
<ID>N_in0</ID>85 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>203</ID>
<type>AA_LABEL</type>
<position>70.5,-62.5</position>
<gparam>LABEL_TEXT S1' S0' Din</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>10</ID>
<type>AA_TOGGLE</type>
<position>24,-3.5</position>
<output>
<ID>OUT_0</ID>4 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>204</ID>
<type>AA_LABEL</type>
<position>70.5,-70.5</position>
<gparam>LABEL_TEXT S1' S0 Din</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>205</ID>
<type>AA_LABEL</type>
<position>71,-78</position>
<gparam>LABEL_TEXT S1 S0' Din</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>12</ID>
<type>AA_LABEL</type>
<position>1,-6.5</position>
<gparam>LABEL_TEXT MUX</gparam>
<gparam>TEXT_HEIGHT 5</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>206</ID>
<type>AA_LABEL</type>
<position>71.5,-86</position>
<gparam>LABEL_TEXT S1 S0 Din</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>207</ID>
<type>AA_LABEL</type>
<position>81.5,-63</position>
<gparam>LABEL_TEXT D0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>14</ID>
<type>AA_LABEL</type>
<position>15,-6.5</position>
<gparam>LABEL_TEXT D0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>208</ID>
<type>AA_LABEL</type>
<position>81.5,-71</position>
<gparam>LABEL_TEXT D1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>15</ID>
<type>AA_LABEL</type>
<position>17.5,-9</position>
<gparam>LABEL_TEXT D1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>209</ID>
<type>AA_LABEL</type>
<position>81.5,-79</position>
<gparam>LABEL_TEXT D2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>210</ID>
<type>AA_LABEL</type>
<position>81.5,-87</position>
<gparam>LABEL_TEXT D3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>17</ID>
<type>AA_LABEL</type>
<position>24,-1</position>
<gparam>LABEL_TEXT S0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>211</ID>
<type>AA_LABEL</type>
<position>61,-52.5</position>
<gparam>LABEL_TEXT 1 X 4 De-mux</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>19</ID>
<type>AE_MUX_4x1</type>
<position>49,-8</position>
<input>
<ID>IN_0</ID>7 </input>
<input>
<ID>IN_1</ID>6 </input>
<input>
<ID>IN_2</ID>5 </input>
<input>
<ID>IN_3</ID>10 </input>
<output>
<ID>OUT</ID>13 </output>
<input>
<ID>SEL_0</ID>9 </input>
<input>
<ID>SEL_1</ID>8 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>21</ID>
<type>AA_TOGGLE</type>
<position>38,-5</position>
<output>
<ID>OUT_0</ID>10 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>23</ID>
<type>AA_TOGGLE</type>
<position>44,-7</position>
<output>
<ID>OUT_0</ID>5 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>25</ID>
<type>AA_TOGGLE</type>
<position>38,-9</position>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>27</ID>
<type>AA_TOGGLE</type>
<position>43.5,-11</position>
<output>
<ID>OUT_0</ID>7 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>29</ID>
<type>AA_TOGGLE</type>
<position>46,0</position>
<output>
<ID>OUT_0</ID>8 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>31</ID>
<type>AA_TOGGLE</type>
<position>52.5,0</position>
<output>
<ID>OUT_0</ID>9 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>33</ID>
<type>GA_LED</type>
<position>53,-8</position>
<input>
<ID>N_in0</ID>13 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>34</ID>
<type>AA_LABEL</type>
<position>41,-11</position>
<gparam>LABEL_TEXT D0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>35</ID>
<type>AA_LABEL</type>
<position>35,-8.5</position>
<gparam>LABEL_TEXT D1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>36</ID>
<type>AA_LABEL</type>
<position>41,-6.5</position>
<gparam>LABEL_TEXT D2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>37</ID>
<type>AA_LABEL</type>
<position>35.5,-4.5</position>
<gparam>LABEL_TEXT D3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>38</ID>
<type>AA_LABEL</type>
<position>45.5,2.5</position>
<gparam>LABEL_TEXT S0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>40</ID>
<type>AI_MUX_8x1</type>
<position>79,-8</position>
<input>
<ID>IN_0</ID>20 </input>
<input>
<ID>IN_1</ID>21 </input>
<input>
<ID>IN_2</ID>22 </input>
<input>
<ID>IN_3</ID>23 </input>
<input>
<ID>IN_4</ID>27 </input>
<input>
<ID>IN_5</ID>26 </input>
<input>
<ID>IN_6</ID>25 </input>
<input>
<ID>IN_7</ID>17 </input>
<output>
<ID>OUT</ID>69 </output>
<input>
<ID>SEL_0</ID>29 </input>
<input>
<ID>SEL_1</ID>28 </input>
<input>
<ID>SEL_2</ID>30 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>42</ID>
<type>AA_TOGGLE</type>
<position>66.5,-1.5</position>
<output>
<ID>OUT_0</ID>25 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>44</ID>
<type>AA_TOGGLE</type>
<position>66.5,-4</position>
<output>
<ID>OUT_0</ID>26 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>46</ID>
<type>AA_TOGGLE</type>
<position>66.5,-9</position>
<output>
<ID>OUT_0</ID>23 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>48</ID>
<type>AA_TOGGLE</type>
<position>66.5,-11.5</position>
<output>
<ID>OUT_0</ID>22 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>50</ID>
<type>AA_TOGGLE</type>
<position>66.5,-14</position>
<output>
<ID>OUT_0</ID>21 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>51</ID>
<type>AA_TOGGLE</type>
<position>66.5,-16.5</position>
<output>
<ID>OUT_0</ID>20 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>52</ID>
<type>AA_TOGGLE</type>
<position>66.5,1</position>
<output>
<ID>OUT_0</ID>17 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>53</ID>
<type>AA_TOGGLE</type>
<position>66.5,-6.5</position>
<output>
<ID>OUT_0</ID>27 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>54</ID>
<type>AA_TOGGLE</type>
<position>77.5,2.5</position>
<output>
<ID>OUT_0</ID>30 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>55</ID>
<type>AA_TOGGLE</type>
<position>80.5,2.5</position>
<output>
<ID>OUT_0</ID>28 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>56</ID>
<type>AA_TOGGLE</type>
<position>83.5,2.5</position>
<output>
<ID>OUT_0</ID>29 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>57</ID>
<type>GA_LED</type>
<position>83,-8</position>
<input>
<ID>N_in0</ID>69 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>58</ID>
<type>AA_LABEL</type>
<position>63.5,-8.5</position>
<gparam>LABEL_TEXT D3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>59</ID>
<type>AA_LABEL</type>
<position>63.5,-11</position>
<gparam>LABEL_TEXT D2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>60</ID>
<type>AA_LABEL</type>
<position>63.5,-13.5</position>
<gparam>LABEL_TEXT D1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>61</ID>
<type>AA_LABEL</type>
<position>63.5,-16</position>
<gparam>LABEL_TEXT D0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>62</ID>
<type>AA_LABEL</type>
<position>63.5,-6</position>
<gparam>LABEL_TEXT D4</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>63</ID>
<type>AA_LABEL</type>
<position>63.5,-3.5</position>
<gparam>LABEL_TEXT D5</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>64</ID>
<type>AA_LABEL</type>
<position>63.5,-1</position>
<gparam>LABEL_TEXT D6</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>65</ID>
<type>AA_LABEL</type>
<position>63.5,1.5</position>
<gparam>LABEL_TEXT D7</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>66</ID>
<type>AA_LABEL</type>
<position>52.5,2.5</position>
<gparam>LABEL_TEXT S1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>67</ID>
<type>AA_LABEL</type>
<position>77.5,5</position>
<gparam>LABEL_TEXT S0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>68</ID>
<type>AA_LABEL</type>
<position>80.5,5</position>
<gparam>LABEL_TEXT S1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>69</ID>
<type>AA_LABEL</type>
<position>83.5,5</position>
<gparam>LABEL_TEXT S2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>70</ID>
<type>AA_LABEL</type>
<position>2,-63.5</position>
<gparam>LABEL_TEXT DE-MUX</gparam>
<gparam>TEXT_HEIGHT 8</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>105</ID>
<type>AA_LABEL</type>
<position>21.5,4</position>
<gparam>LABEL_TEXT 2 X 1 mux</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>107</ID>
<type>AA_LABEL</type>
<position>48,5.5</position>
<gparam>LABEL_TEXT 4 X 1 mux</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>108</ID>
<type>AA_LABEL</type>
<position>74,8.5</position>
<gparam>LABEL_TEXT 8 X 1 mux</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>114</ID>
<type>AA_TOGGLE</type>
<position>114,-31.5</position>
<output>
<ID>OUT_0</ID>57 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>115</ID>
<type>AA_TOGGLE</type>
<position>123,-31.5</position>
<output>
<ID>OUT_0</ID>56 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>116</ID>
<type>AA_TOGGLE</type>
<position>131,-31.5</position>
<output>
<ID>OUT_0</ID>52 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>117</ID>
<type>AE_SMALL_INVERTER</type>
<position>118,-35.5</position>
<input>
<ID>IN_0</ID>57 </input>
<output>
<ID>OUT_0</ID>54 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>118</ID>
<type>AE_SMALL_INVERTER</type>
<position>127,-35.5</position>
<input>
<ID>IN_0</ID>56 </input>
<output>
<ID>OUT_0</ID>53 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>123</ID>
<type>AA_LABEL</type>
<position>123,-28.5</position>
<gparam>LABEL_TEXT S0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>124</ID>
<type>AA_LABEL</type>
<position>114,-28.5</position>
<gparam>LABEL_TEXT S1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>125</ID>
<type>AA_LABEL</type>
<position>131,-28.5</position>
<gparam>LABEL_TEXT Din</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>126</ID>
<type>GA_LED</type>
<position>159,-43.5</position>
<input>
<ID>N_in0</ID>64 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>127</ID>
<type>GA_LED</type>
<position>159.5,-53.5</position>
<input>
<ID>N_in0</ID>61 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>128</ID>
<type>GA_LED</type>
<position>160,-63.5</position>
<input>
<ID>N_in0</ID>62 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>129</ID>
<type>GA_LED</type>
<position>160,-73</position>
<input>
<ID>N_in0</ID>63 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>134</ID>
<type>AA_LABEL</type>
<position>164.5,-43</position>
<gparam>LABEL_TEXT D0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>135</ID>
<type>AA_LABEL</type>
<position>165,-53</position>
<gparam>LABEL_TEXT D1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>136</ID>
<type>AA_LABEL</type>
<position>165,-63</position>
<gparam>LABEL_TEXT D2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>137</ID>
<type>AA_LABEL</type>
<position>165,-72.5</position>
<gparam>LABEL_TEXT D3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>138</ID>
<type>AA_TOGGLE</type>
<position>104,-31.5</position>
<output>
<ID>OUT_0</ID>60 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>139</ID>
<type>AE_SMALL_INVERTER</type>
<position>108.5,-35.5</position>
<input>
<ID>IN_0</ID>60 </input>
<output>
<ID>OUT_0</ID>55 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>141</ID>
<type>AA_AND4</type>
<position>155,-43.5</position>
<input>
<ID>IN_0</ID>53 </input>
<input>
<ID>IN_1</ID>54 </input>
<input>
<ID>IN_2</ID>55 </input>
<input>
<ID>IN_3</ID>52 </input>
<output>
<ID>OUT</ID>64 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>142</ID>
<type>AA_AND4</type>
<position>155.5,-53.5</position>
<input>
<ID>IN_0</ID>56 </input>
<input>
<ID>IN_1</ID>54 </input>
<input>
<ID>IN_2</ID>55 </input>
<input>
<ID>IN_3</ID>52 </input>
<output>
<ID>OUT</ID>61 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>143</ID>
<type>AA_AND4</type>
<position>156,-63.5</position>
<input>
<ID>IN_0</ID>53 </input>
<input>
<ID>IN_1</ID>57 </input>
<input>
<ID>IN_2</ID>55 </input>
<input>
<ID>IN_3</ID>52 </input>
<output>
<ID>OUT</ID>62 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>144</ID>
<type>AA_AND4</type>
<position>156,-73</position>
<input>
<ID>IN_0</ID>56 </input>
<input>
<ID>IN_1</ID>57 </input>
<input>
<ID>IN_2</ID>55 </input>
<input>
<ID>IN_3</ID>52 </input>
<output>
<ID>OUT</ID>63 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>146</ID>
<type>AA_AND4</type>
<position>156,-92</position>
<input>
<ID>IN_0</ID>56 </input>
<input>
<ID>IN_1</ID>54 </input>
<input>
<ID>IN_2</ID>60 </input>
<input>
<ID>IN_3</ID>52 </input>
<output>
<ID>OUT</ID>66 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>147</ID>
<type>AA_AND4</type>
<position>156,-101.5</position>
<input>
<ID>IN_0</ID>53 </input>
<input>
<ID>IN_1</ID>57 </input>
<input>
<ID>IN_2</ID>60 </input>
<input>
<ID>IN_3</ID>52 </input>
<output>
<ID>OUT</ID>67 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>148</ID>
<type>AA_AND4</type>
<position>156,-111</position>
<input>
<ID>IN_0</ID>56 </input>
<input>
<ID>IN_1</ID>57 </input>
<input>
<ID>IN_2</ID>60 </input>
<input>
<ID>IN_3</ID>52 </input>
<output>
<ID>OUT</ID>68 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>149</ID>
<type>AA_AND4</type>
<position>156,-82.5</position>
<input>
<ID>IN_0</ID>53 </input>
<input>
<ID>IN_1</ID>54 </input>
<input>
<ID>IN_2</ID>60 </input>
<input>
<ID>IN_3</ID>52 </input>
<output>
<ID>OUT</ID>65 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>150</ID>
<type>GA_LED</type>
<position>160,-82.5</position>
<input>
<ID>N_in0</ID>65 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>151</ID>
<type>GA_LED</type>
<position>160,-92</position>
<input>
<ID>N_in0</ID>66 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>152</ID>
<type>GA_LED</type>
<position>160,-101.5</position>
<input>
<ID>N_in0</ID>67 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>153</ID>
<type>GA_LED</type>
<position>160,-111</position>
<input>
<ID>N_in0</ID>68 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>155</ID>
<type>AA_LABEL</type>
<position>165,-82</position>
<gparam>LABEL_TEXT D4</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>156</ID>
<type>AA_LABEL</type>
<position>165,-91.5</position>
<gparam>LABEL_TEXT D5</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>157</ID>
<type>AA_LABEL</type>
<position>165.5,-101</position>
<gparam>LABEL_TEXT D6</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>158</ID>
<type>AA_LABEL</type>
<position>165.5,-110</position>
<gparam>LABEL_TEXT D7</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>160</ID>
<type>AA_LABEL</type>
<position>145,-35.5</position>
<gparam>LABEL_TEXT 1 X 8 De-mux</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>161</ID>
<type>AA_LABEL</type>
<position>104,-28.5</position>
<gparam>LABEL_TEXT S2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>187</ID>
<type>AA_TOGGLE</type>
<position>26.5,-53</position>
<output>
<ID>OUT_0</ID>81 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>188</ID>
<type>AA_TOGGLE</type>
<position>35.5,-53</position>
<output>
<ID>OUT_0</ID>83 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>189</ID>
<type>AA_TOGGLE</type>
<position>43.5,-53</position>
<output>
<ID>OUT_0</ID>79 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>190</ID>
<type>AE_SMALL_INVERTER</type>
<position>30.5,-57</position>
<input>
<ID>IN_0</ID>81 </input>
<output>
<ID>OUT_0</ID>80 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>191</ID>
<type>AE_SMALL_INVERTER</type>
<position>39.5,-57</position>
<input>
<ID>IN_0</ID>83 </input>
<output>
<ID>OUT_0</ID>82 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>192</ID>
<type>AA_AND3</type>
<position>64,-63.5</position>
<input>
<ID>IN_0</ID>80 </input>
<input>
<ID>IN_1</ID>82 </input>
<input>
<ID>IN_2</ID>79 </input>
<output>
<ID>OUT</ID>86 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<wire>
<ID>1</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19.5,-7,22,-7</points>
<connection>
<GID>2</GID>
<name>IN_1</name></connection>
<connection>
<GID>4</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22,-9,22,-9</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26,-8,26,-8</points>
<connection>
<GID>2</GID>
<name>OUT</name></connection>
<connection>
<GID>8</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24,-5.5,24,-5.5</points>
<connection>
<GID>2</GID>
<name>SEL_0</name></connection>
<connection>
<GID>10</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>46,-7,46,-7</points>
<connection>
<GID>23</GID>
<name>OUT_0</name></connection>
<connection>
<GID>19</GID>
<name>IN_2</name></connection></vsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>40,-9,46,-9</points>
<connection>
<GID>19</GID>
<name>IN_1</name></connection>
<connection>
<GID>25</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45.5,-11,46,-11</points>
<connection>
<GID>19</GID>
<name>IN_0</name></connection>
<connection>
<GID>27</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>46,-3,46,-2</points>
<connection>
<GID>29</GID>
<name>OUT_0</name></connection>
<intersection>-3 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>46,-3,49,-3</points>
<connection>
<GID>19</GID>
<name>SEL_1</name></connection>
<intersection>46 0</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52.5,-3,52.5,-2</points>
<connection>
<GID>31</GID>
<name>OUT_0</name></connection>
<intersection>-3 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50,-3,52.5,-3</points>
<connection>
<GID>19</GID>
<name>SEL_0</name></connection>
<intersection>52.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>40,-5,46,-5</points>
<connection>
<GID>19</GID>
<name>IN_3</name></connection>
<connection>
<GID>21</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52,-8,52,-8</points>
<connection>
<GID>33</GID>
<name>N_in0</name></connection>
<connection>
<GID>19</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>68.5,1,76,1</points>
<connection>
<GID>52</GID>
<name>OUT_0</name></connection>
<intersection>76 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>76,-4.5,76,1</points>
<connection>
<GID>40</GID>
<name>IN_7</name></connection>
<intersection>1 1</intersection></vsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>68.5,-16.5,76,-16.5</points>
<connection>
<GID>51</GID>
<name>OUT_0</name></connection>
<intersection>76 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>76,-16.5,76,-11.5</points>
<connection>
<GID>40</GID>
<name>IN_0</name></connection>
<intersection>-16.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>72,-14,72,-10.5</points>
<intersection>-14 1</intersection>
<intersection>-10.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>68.5,-14,72,-14</points>
<connection>
<GID>50</GID>
<name>OUT_0</name></connection>
<intersection>72 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>72,-10.5,76,-10.5</points>
<connection>
<GID>40</GID>
<name>IN_1</name></connection>
<intersection>72 0</intersection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>68.5,-11.5,71,-11.5</points>
<connection>
<GID>48</GID>
<name>OUT_0</name></connection>
<intersection>71 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>71,-11.5,71,-9.5</points>
<intersection>-11.5 1</intersection>
<intersection>-9.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>71,-9.5,76,-9.5</points>
<connection>
<GID>40</GID>
<name>IN_2</name></connection>
<intersection>71 3</intersection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>72,-9,72,-8.5</points>
<intersection>-9 1</intersection>
<intersection>-8.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>68.5,-9,72,-9</points>
<connection>
<GID>46</GID>
<name>OUT_0</name></connection>
<intersection>72 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>72,-8.5,76,-8.5</points>
<connection>
<GID>40</GID>
<name>IN_3</name></connection>
<intersection>72 0</intersection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73.5,-5.5,73.5,-1.5</points>
<intersection>-5.5 2</intersection>
<intersection>-1.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>68.5,-1.5,73.5,-1.5</points>
<connection>
<GID>42</GID>
<name>OUT_0</name></connection>
<intersection>73.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>73.5,-5.5,76,-5.5</points>
<connection>
<GID>40</GID>
<name>IN_6</name></connection>
<intersection>73.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>72.5,-6.5,72.5,-4</points>
<intersection>-6.5 2</intersection>
<intersection>-4 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>68.5,-4,72.5,-4</points>
<connection>
<GID>44</GID>
<name>OUT_0</name></connection>
<intersection>72.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>72.5,-6.5,76,-6.5</points>
<connection>
<GID>40</GID>
<name>IN_5</name></connection>
<intersection>72.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>72,-7.5,72,-6.5</points>
<intersection>-7.5 2</intersection>
<intersection>-6.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>68.5,-6.5,72,-6.5</points>
<connection>
<GID>53</GID>
<name>OUT_0</name></connection>
<intersection>72 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>72,-7.5,76,-7.5</points>
<connection>
<GID>40</GID>
<name>IN_4</name></connection>
<intersection>72 0</intersection></hsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80.5,-1,80.5,0.5</points>
<connection>
<GID>55</GID>
<name>OUT_0</name></connection>
<intersection>-1 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>79,-2.5,79,-1</points>
<connection>
<GID>40</GID>
<name>SEL_1</name></connection>
<intersection>-1 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>79,-1,80.5,-1</points>
<intersection>79 1</intersection>
<intersection>80.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>83.5,-1.5,83.5,0.5</points>
<connection>
<GID>56</GID>
<name>OUT_0</name></connection>
<intersection>-1.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>80,-2.5,80,-1.5</points>
<connection>
<GID>40</GID>
<name>SEL_0</name></connection>
<intersection>-1.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>80,-1.5,83.5,-1.5</points>
<intersection>80 1</intersection>
<intersection>83.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>77.5,-1,77.5,0.5</points>
<connection>
<GID>54</GID>
<name>OUT_0</name></connection>
<intersection>-1 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>78,-2.5,78,-1</points>
<connection>
<GID>40</GID>
<name>SEL_2</name></connection>
<intersection>-1 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>77.5,-1,78,-1</points>
<intersection>77.5 0</intersection>
<intersection>78 1</intersection></hsegment></shape></wire>
<wire>
<ID>52</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>131,-114,131,-33.5</points>
<connection>
<GID>116</GID>
<name>OUT_0</name></connection>
<intersection>-114 5</intersection>
<intersection>-104.5 15</intersection>
<intersection>-95 13</intersection>
<intersection>-85.5 17</intersection>
<intersection>-76 9</intersection>
<intersection>-66.5 7</intersection>
<intersection>-56.5 3</intersection>
<intersection>-46.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>131,-46.5,152,-46.5</points>
<connection>
<GID>141</GID>
<name>IN_3</name></connection>
<intersection>131 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>131,-56.5,152.5,-56.5</points>
<connection>
<GID>142</GID>
<name>IN_3</name></connection>
<intersection>131 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>131,-114,153,-114</points>
<connection>
<GID>148</GID>
<name>IN_3</name></connection>
<intersection>131 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>131,-66.5,153,-66.5</points>
<connection>
<GID>143</GID>
<name>IN_3</name></connection>
<intersection>131 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>131,-76,153,-76</points>
<connection>
<GID>144</GID>
<name>IN_3</name></connection>
<intersection>131 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>131,-95,153,-95</points>
<connection>
<GID>146</GID>
<name>IN_3</name></connection>
<intersection>131 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>131,-104.5,153,-104.5</points>
<connection>
<GID>147</GID>
<name>IN_3</name></connection>
<intersection>131 0</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>131,-85.5,153,-85.5</points>
<connection>
<GID>149</GID>
<name>IN_3</name></connection>
<intersection>131 0</intersection></hsegment></shape></wire>
<wire>
<ID>53</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>127,-98.5,127,-37.5</points>
<connection>
<GID>118</GID>
<name>OUT_0</name></connection>
<intersection>-98.5 7</intersection>
<intersection>-79.5 5</intersection>
<intersection>-60.5 3</intersection>
<intersection>-40.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>127,-40.5,152,-40.5</points>
<connection>
<GID>141</GID>
<name>IN_0</name></connection>
<intersection>127 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>127,-60.5,153,-60.5</points>
<connection>
<GID>143</GID>
<name>IN_0</name></connection>
<intersection>127 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>127,-79.5,153,-79.5</points>
<connection>
<GID>149</GID>
<name>IN_0</name></connection>
<intersection>127 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>127,-98.5,153,-98.5</points>
<connection>
<GID>147</GID>
<name>IN_0</name></connection>
<intersection>127 0</intersection></hsegment></shape></wire>
<wire>
<ID>54</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>117.5,-91,117.5,-37.5</points>
<intersection>-91 7</intersection>
<intersection>-81.5 5</intersection>
<intersection>-52.5 3</intersection>
<intersection>-42.5 1</intersection>
<intersection>-37.5 8</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>117.5,-42.5,152,-42.5</points>
<connection>
<GID>141</GID>
<name>IN_1</name></connection>
<intersection>117.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>117.5,-52.5,152.5,-52.5</points>
<connection>
<GID>142</GID>
<name>IN_1</name></connection>
<intersection>117.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>117.5,-81.5,153,-81.5</points>
<connection>
<GID>149</GID>
<name>IN_1</name></connection>
<intersection>117.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>117.5,-91,153,-91</points>
<connection>
<GID>146</GID>
<name>IN_1</name></connection>
<intersection>117.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>117.5,-37.5,118,-37.5</points>
<connection>
<GID>117</GID>
<name>OUT_0</name></connection>
<intersection>117.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>55</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>108.5,-74,108.5,-37.5</points>
<connection>
<GID>139</GID>
<name>OUT_0</name></connection>
<intersection>-74 7</intersection>
<intersection>-64.5 5</intersection>
<intersection>-54.5 3</intersection>
<intersection>-44.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>108.5,-44.5,152,-44.5</points>
<connection>
<GID>141</GID>
<name>IN_2</name></connection>
<intersection>108.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>108.5,-54.5,152.5,-54.5</points>
<connection>
<GID>142</GID>
<name>IN_2</name></connection>
<intersection>108.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>108.5,-64.5,153,-64.5</points>
<connection>
<GID>143</GID>
<name>IN_2</name></connection>
<intersection>108.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>108.5,-74,153,-74</points>
<connection>
<GID>144</GID>
<name>IN_2</name></connection>
<intersection>108.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>56</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>123,-108,123,-33.5</points>
<connection>
<GID>115</GID>
<name>OUT_0</name></connection>
<intersection>-108 11</intersection>
<intersection>-89 9</intersection>
<intersection>-70 3</intersection>
<intersection>-50.5 1</intersection>
<intersection>-33.5 12</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>123,-50.5,152.5,-50.5</points>
<connection>
<GID>142</GID>
<name>IN_0</name></connection>
<intersection>123 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>123,-70,153,-70</points>
<connection>
<GID>144</GID>
<name>IN_0</name></connection>
<intersection>123 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>123,-89,153,-89</points>
<connection>
<GID>146</GID>
<name>IN_0</name></connection>
<intersection>123 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>123,-108,153,-108</points>
<connection>
<GID>148</GID>
<name>IN_0</name></connection>
<intersection>123 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>123,-33.5,127,-33.5</points>
<connection>
<GID>118</GID>
<name>IN_0</name></connection>
<intersection>123 0</intersection></hsegment></shape></wire>
<wire>
<ID>57</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>114,-110,114,-33.5</points>
<connection>
<GID>114</GID>
<name>OUT_0</name></connection>
<intersection>-110 9</intersection>
<intersection>-100.5 7</intersection>
<intersection>-72 3</intersection>
<intersection>-62.5 1</intersection>
<intersection>-33.5 10</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>114,-62.5,153,-62.5</points>
<connection>
<GID>143</GID>
<name>IN_1</name></connection>
<intersection>114 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>114,-72,153,-72</points>
<connection>
<GID>144</GID>
<name>IN_1</name></connection>
<intersection>114 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>114,-100.5,153,-100.5</points>
<connection>
<GID>147</GID>
<name>IN_1</name></connection>
<intersection>114 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>114,-110,153,-110</points>
<connection>
<GID>148</GID>
<name>IN_1</name></connection>
<intersection>114 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>114,-33.5,118,-33.5</points>
<connection>
<GID>117</GID>
<name>IN_0</name></connection>
<intersection>114 0</intersection></hsegment></shape></wire>
<wire>
<ID>60</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>104,-112,104,-33.5</points>
<connection>
<GID>138</GID>
<name>OUT_0</name></connection>
<intersection>-112 5</intersection>
<intersection>-102.5 7</intersection>
<intersection>-93 3</intersection>
<intersection>-83.5 1</intersection>
<intersection>-33.5 8</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>104,-83.5,153,-83.5</points>
<connection>
<GID>149</GID>
<name>IN_2</name></connection>
<intersection>104 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>104,-93,153,-93</points>
<connection>
<GID>146</GID>
<name>IN_2</name></connection>
<intersection>104 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>104,-112,153,-112</points>
<connection>
<GID>148</GID>
<name>IN_2</name></connection>
<intersection>104 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>104,-102.5,153,-102.5</points>
<connection>
<GID>147</GID>
<name>IN_2</name></connection>
<intersection>104 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>104,-33.5,108.5,-33.5</points>
<connection>
<GID>139</GID>
<name>IN_0</name></connection>
<intersection>104 0</intersection></hsegment></shape></wire>
<wire>
<ID>61</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>158.5,-53.5,158.5,-53.5</points>
<connection>
<GID>127</GID>
<name>N_in0</name></connection>
<connection>
<GID>142</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>62</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>159,-63.5,159,-63.5</points>
<connection>
<GID>128</GID>
<name>N_in0</name></connection>
<connection>
<GID>143</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>63</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>159,-73,159,-73</points>
<connection>
<GID>129</GID>
<name>N_in0</name></connection>
<connection>
<GID>144</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>64</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>158,-43.5,158,-43.5</points>
<connection>
<GID>126</GID>
<name>N_in0</name></connection>
<connection>
<GID>141</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>65</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>159,-82.5,159,-82.5</points>
<connection>
<GID>149</GID>
<name>OUT</name></connection>
<connection>
<GID>150</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>66</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>159,-92,159,-92</points>
<connection>
<GID>146</GID>
<name>OUT</name></connection>
<connection>
<GID>151</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>67</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>159,-101.5,159,-101.5</points>
<connection>
<GID>147</GID>
<name>OUT</name></connection>
<connection>
<GID>152</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>68</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>159,-111,159,-111</points>
<connection>
<GID>148</GID>
<name>OUT</name></connection>
<connection>
<GID>153</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>69</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>82,-8,82,-8</points>
<connection>
<GID>40</GID>
<name>OUT</name></connection>
<connection>
<GID>57</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>79</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>43.5,-89.5,43.5,-55</points>
<connection>
<GID>189</GID>
<name>OUT_0</name></connection>
<intersection>-89.5 7</intersection>
<intersection>-81.5 5</intersection>
<intersection>-73.5 3</intersection>
<intersection>-65.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>43.5,-65.5,61,-65.5</points>
<connection>
<GID>192</GID>
<name>IN_2</name></connection>
<intersection>43.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>43.5,-73.5,61,-73.5</points>
<connection>
<GID>193</GID>
<name>IN_2</name></connection>
<intersection>43.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>43.5,-81.5,61,-81.5</points>
<connection>
<GID>194</GID>
<name>IN_2</name></connection>
<intersection>43.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>43.5,-89.5,61,-89.5</points>
<connection>
<GID>195</GID>
<name>IN_2</name></connection>
<intersection>43.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>80</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30.5,-69.5,30.5,-59</points>
<connection>
<GID>190</GID>
<name>OUT_0</name></connection>
<intersection>-69.5 3</intersection>
<intersection>-61.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30.5,-61.5,61,-61.5</points>
<connection>
<GID>192</GID>
<name>IN_0</name></connection>
<intersection>30.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>30.5,-69.5,61,-69.5</points>
<connection>
<GID>193</GID>
<name>IN_0</name></connection>
<intersection>30.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>81</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26.5,-85.5,26.5,-55</points>
<connection>
<GID>187</GID>
<name>OUT_0</name></connection>
<intersection>-85.5 3</intersection>
<intersection>-77.5 1</intersection>
<intersection>-55 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26.5,-77.5,61,-77.5</points>
<connection>
<GID>194</GID>
<name>IN_0</name></connection>
<intersection>26.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>26.5,-85.5,61,-85.5</points>
<connection>
<GID>195</GID>
<name>IN_0</name></connection>
<intersection>26.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>26.5,-55,30.5,-55</points>
<connection>
<GID>190</GID>
<name>IN_0</name></connection>
<intersection>26.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>82</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39.5,-79.5,39.5,-59</points>
<connection>
<GID>191</GID>
<name>OUT_0</name></connection>
<intersection>-79.5 3</intersection>
<intersection>-63.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>39.5,-63.5,61,-63.5</points>
<connection>
<GID>192</GID>
<name>IN_1</name></connection>
<intersection>39.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>39.5,-79.5,61,-79.5</points>
<connection>
<GID>194</GID>
<name>IN_1</name></connection>
<intersection>39.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>83</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35.5,-87.5,35.5,-55</points>
<connection>
<GID>188</GID>
<name>OUT_0</name></connection>
<intersection>-87.5 3</intersection>
<intersection>-71.5 1</intersection>
<intersection>-55 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35.5,-71.5,61,-71.5</points>
<connection>
<GID>193</GID>
<name>IN_1</name></connection>
<intersection>35.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>35.5,-87.5,61,-87.5</points>
<connection>
<GID>195</GID>
<name>IN_1</name></connection>
<intersection>35.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>35.5,-55,39.5,-55</points>
<connection>
<GID>191</GID>
<name>IN_0</name></connection>
<intersection>35.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>84</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>67,-79.5,76,-79.5</points>
<connection>
<GID>194</GID>
<name>OUT</name></connection>
<connection>
<GID>201</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>85</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>67,-87.5,76,-87.5</points>
<connection>
<GID>195</GID>
<name>OUT</name></connection>
<connection>
<GID>202</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>86</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>67,-63.5,75.5,-63.5</points>
<connection>
<GID>192</GID>
<name>OUT</name></connection>
<connection>
<GID>199</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>87</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>67,-71.5,75.5,-71.5</points>
<connection>
<GID>193</GID>
<name>OUT</name></connection>
<connection>
<GID>200</GID>
<name>N_in0</name></connection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,0,145.8,-73.7</PageViewport></page 1>
<page 2>
<PageViewport>0,0,145.8,-73.7</PageViewport></page 2>
<page 3>
<PageViewport>0,0,145.8,-73.7</PageViewport></page 3>
<page 4>
<PageViewport>0,0,145.8,-73.7</PageViewport></page 4>
<page 5>
<PageViewport>0,0,145.8,-73.7</PageViewport></page 5>
<page 6>
<PageViewport>0,0,145.8,-73.7</PageViewport></page 6>
<page 7>
<PageViewport>0,0,145.8,-73.7</PageViewport></page 7>
<page 8>
<PageViewport>0,0,145.8,-73.7</PageViewport></page 8>
<page 9>
<PageViewport>0,0,145.8,-73.7</PageViewport></page 9></circuit>